Entity evbx1_ep2m_tb is
End evbx1_ep2m_tb;
