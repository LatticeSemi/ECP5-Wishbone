`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2021.04.107"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
KS4j+re0KO85GJkuS0W+2MR6VFpwVGCEBzrnnCFDcPU6x0lNgfF5qQNs3fsEqpHVvzlg9WYXcRa/
Y6hQAAADgKVnzRrD33n2DN+PV+sSuw3knmwU5zLlSD+Jt6W2g7b55jszmBatbaV3LJQi0QCdRbPt
eHsrwFVBavZT2ttswLnwx+elT/MNF0Fb0rgosjMHhDWF0ASx8cm3LAVxIqLVebrwNf4xl2Jwo7KQ
n0D9+LIEOIU93hC+aeulAtfDjq5E+f0NfMHkHh78zfLQ0kEby6KlMYee5AF53vvJ5ERmlF3RUbLz
ty5JRUm2yGV1WfER5uBlhHCF19Im9h9MHuzsv+==
`protect key_keyowner= "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-3", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 128)
`protect key_block
aDXC881+wcKu7aMeU8cGTFcDVWrZYOuaCUI2ZXnztnA4TMdGc0CIWuOuo7woLbo1d8zzggIRQVTc
/qAH7hMOh7SU2y/ObfU3RO4AiC0P6sQYn5QfWrHeNigBulFLD4FcvOSs78Yy7w75LP/K/xu3tETI
8Qv4E8CBuBmErcz1ZW/=

`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 642592)
`protect data_block
away4wqJ0ZObdLfFSDKe0NffzHpasfWcx1MOZ/C9p0+YQM1OJ35mgXROUpoKmTjNDjaXysXQdQmy
ZCH4w3QXvmYla+iWqyNiMvT/N0llL3QiRKiUE8oYPjiRQjX1SMRxsGn1fubcAXGEpofzNg+F+PGA
PpLTmi0Mm93SDxBud0aFu0ohXAg1HY3b1nOeKUhfcY5AFaZJaIKzMrOcbZ18+VNuaeyarwVz//4M
Y+G2HL7xm4Xk/xvAq13maPf+UUeDrd7lpFIj2JzBZ5z3SnblYYJXD0fhnwxkC+Nfuzf5KGmgPcs3
RGRLpiNR+bLBhTJb9dGY4qNLzjpHNBdH++izEboRkSS8YKuhzxCW3/oTDHlA7kkZaLqDUQnD/j9o
G85e+CHSPHyPmvSPGECb4eY9LwfdN7YlE9m62rfDRhC673MlgqXuTuUT3LRzFd9Znn627NbrQxx5
qyzqRKm0/h9b2TU7GR+t0IfMfxbzNBxmzJz4TPGBZbs0Ss3I2qJcUdK24LC/lc3enCG1h8Bi9BPg
jCVi92dQgB6Bsh6dsYOl1/6mysZT6PuQnmgCrxzG0AwAC6OZEbVBKr7e6X5X7t2p6ZsDAxwR4omp
e6LKU28swyHvonV8+DFJeURvOsS1znvR2ZJozJOXePrUZgrhENmzWQHwvW+JOGZ9X26SRmGhPysQ
YQCALXFOyOObAxVq3Mp57JaGPDaslzKjfAeOO4hOfAR8Uq7+mGvLbXjIfu8BesejZ51kn9zhE1bq
UL9zf6g57wyvnnS+KJ/hOrOugsYjFAuJFC15GyPQVkOFhFUiYy81FKg8QzLskBbyxxF80y/THuiy
D7d7MXy8VftQBOqT8seESZKqhkUxeQKYN52OMzEPOtunJhHkLbFlU7oUe8j0fxlCZXwncHKcPHC3
AnUoJXUgI+KyErJ/z5GS6I77kOTOCRju83n16Hi7pA5Tq0VT+1d3MyTgLqljiR3cm9g2HqZm1k3O
5cslqyutRfSuBY54muPITHDpSzR4uR5yBoj99QhYLZQ9n222Ua5vU0BF/RM1oy/iCp/xQs1t369v
GM5A+fUIhmKBYgSA6gi0l8y6/brIU7QVN/97BRgn3Dd4dEW/mOrdMgZnlse3AIen9TCCyLw/LfBD
dbantit8UJePjDQvxNril7kU+dhtE99wUmFBRTtly+IebsSdnz1z1yunsng0QYloxpPMB6va6Smh
GTSKe7q30/THchHpjKHRMvBk22t3sUrP39EZodon0sygsVUQIdiFfOTRL/JXF/hR1KhSSthJaKWT
GGH+3m7ukUqtQos7HSjH94WvzBe0cqIFIVWvPPN4AZVSS0za35fKmb8LfUNSr7V4bIyicwedR0Pz
22waPvwLMzYHM0157ZvwDMriMy1mJEfSWwvvSICz5gT8f8iSbpUBkiVXOFh0S2oFmN4z/XieMm6O
K9iY8W26ihjlP57abnoq/kTtXoMVOmmnNkQhFHyI3TsmipYbxLG5openg/wWPJXe3qBbw/GO0Nrz
YVyzQjEzYy5sAIqVfIy1f9pmxLHhyR5pO3z20Ubljfzh24Jv8Q9ySL2JLww4Qx9Ll8lZoLOtvA0F
vQHej/TjuXvW8n2JyryZ1oNcW//EEBHDow71+4p01F+GfLhP5kAr1iWOr+w6zwBZAoeKcby9D8I5
yEUUqIS5YyKwL8uhUgCaSj0tSOVVs85jHBF9sp4+gDsPVHk1vntT4Ld56nQdm+FT0Rp8B08C8sCT
1CargUnGCiWAoPlRJ+RuzRDpYTbA9eAoS2ez3g4DniI8JuvdMx+LPpbKA/M7//4f4rkZ/NSbs/Ik
P9rv9AaTefRhNFx0RyauVZ5xEBaP+AcQ4j6aAXlcHeXzTOz7L5Vn8uEm2HJB72yU39JpT3Q5YvS0
vYx8jfciZI2aLJDDfqrDb8IDHcMSxy6orlXT/VzF16umspAkjq/wecAjWhtPZOTuwx4UcgiA1rF3
RkWdzLqogavm068MJAINzgzzMlFicrlNOEMDD95VCDEpEZNHByZie0yvok4AE3MMu1P/sFQ48OG5
DpOFCAH9DmtPOP/e2wrl+/OiuKnCsvMh12ocGMGtUEx7/n0w5euN3QjCZLw+Fvpm4GsN8JmmeRg9
9SqyCeTXZuYCFzWoRp5idaBO7Jb1lvkUZVxdAwwIUhMLBKHIJiXE4CPPm5Cetoyw8Pxgy5ObPD+8
iaETcnPixyqMQ+sOK3g/HrAGHi6XsfPspSWqWww92DuTuislKlkUuUHqBkwHeLtdZfEbmJAYpbyl
8GB5LyaBRvapSWXzdNDfhzqIuqqojV8o2i4L6bff0Qi+ccI09dMJPPOfJGd1jVHc/U1SQtA/cb1Y
+OeUO2PucvpO+ZjdPJMEEvbI2gV/6UqdFM8uiRXCE5J5jqGgy8NUg+Axzz/AJfJjLSCKW36aqIuY
R7QTV4IMdn+TxO+u+Z/Pcy27sA28MBENfCLAftFB70LMlcFF1g6841mL6XdeGWDu8wHmZy3fjIWB
y1OkCweqHKO5bSvf1r+/kE/YtcQ0t7vyps9yyBZezp6q3yif9VinK8s74IbGyOmH0Z0Mfb6WHyGJ
TtATe2+5Nx627++X6x9O420Sn0FoIdw6D+jZG0assYvfRXn2vJ+IW3IQFvWn3yi/exy20I4gry5c
Vc/O4hGKYBcGakspBfxXCFBdoD4F7XRbYpzeiC/yhyrNTfz4pNEbFPDHn5AxDvEXCqKCn+G3k3cv
Olh1yT9MlWGNs4zunk+VKTCEuMoFUrZHKdsM+7lV849OtAPc32fpexM7M1VpKWR617eaRTuvt/y0
I7dCbeWMxq+nO7WEZnYX5a2up0GsJjsSNSspAgP+KszqyWHRLVc3AmREzhgTPrKFH/zz8r7Tb4M7
Lwhy5l2Ei6EoDizumF7xkkank4669NT3W7CfgpzPA5V1Sl9tZOFJKQ9hjsKw/ecnkE1b3AyOS50/
vFQK8yMsuDt3N+7ImuYaxuBJ8XesY4SQZQqpDn4vdjzbfWl9S3HgP9QRbUtDi2FpTYFBUVFrntF8
S9vyH+8NWp2sfXZx1bDkYEchbBIwyZpCLKQGbD3AcO5DX0u397Lsaxe8MHFQAelqoU6le+/njFKn
WEJW+1G0ampT9X2G4foMubzeWs9K2leCv79yx6jruRgoU1vyylur25g+9+cqdZwiL1q28r1IL+SS
vy008MvI8IWMHnaPh2loXL9n2zYk0j4/5JQPnRhIxR9lyExUsVBMmavoVBqXOTaVSDki0cVF2i5t
77o5rXNfXAc6vLAXhmKipwsSqKt20QD5NVfhms2BhhW0sweIKK9xW5PmRA4/IaHtZoAXZgaYCs3O
O+4YAVMJrC2A6pbKSfUatz+4RX19g87FA3WEp0quAJTWyxKtKknSZCwKpgtQuhOp1kcFE9HyM6zg
XZwG6bo4/tQKR6m8NijLyC95q2x2kFnz6WU0i4bVar2e8baUVZTFpydXaSC1TR6yftBEzZWjfa7n
ZTV5DWX5UdjRrwykLDouP4HFriltuomADa+JClzkPwSlGAAcCmUg9Ya29fGQDEQZPq6T24IB+oAL
qR+N0nUZmr9Y3xQvy8CeD4EfX/VUuL1w/s4K60VO83KRQ3ugbTMOWQccpVQKsgTz60cX9U1GYpDY
+SSi/QlRGIFh3T7EdE0fttIBA+AoFo66z46l6o+lpTilIzHfs+aj2CveHfM62zoyJw2PuG6g7w0S
KTOaN3SRfj8a9FZCL6Bdxsm2mo+6+GDQXvq8lzK8vkpZOY8nJjfzHNt0ZKcTdgmSYh4fxZm/7Sr3
JiHUsgR8VScFh9HG6+H4fM5zwLnjA9Q1jnYRXgGITIxCdMZrsRTWPKDz7Fp4YbiijATUQ0qnpQHD
gvtSi+3jet5tcd8PCsbJq/Q3PmuimyQAjj/zykYlteo0X+6uD23Xcpmig4uCZ7GCmIQpoGL27Gm0
jUlwio7+cg/c+7EMnTSARDdbOFUlc9tFwYfjQLup3VG1Rwvn+naLcL3TEocZiHOeDL9B5SW4Hv7Y
1rBQIKkLLhVIohl3JSiBzPGQ+ClVK21qHSbK/6rmvJqrhiHsawgzDrBJ7brOhJFdc+gpi5d9orn7
EhfCxUSg3Ndw9zBt329EE/BUTF79pmu+1cB6RnWryZOAyseFsJNtegmCSo3tmdRoVnGFI65R+6cR
0ITzJJKuquR/6xk2bb8bW6xRsFPNX/M39ipugB0s+73XPwnd7NaZ69Qmr8wHhqVOaxS4UA2WS1tD
B1E4x/sFb4wQBE5HWkq6kxpjqFMP9WSUO1reJA2wsyI3dTEHcIbt79Vu/anfEifDa5m8afx5ed+c
5n+CJ/ptxhGUd6vU4AizqHgjs/oer6rfq1LZXlDAdhoU1Rj9YxaZmsguE2bMFp9oAZx18ohsnJaY
7xCAu86vykX2bAHZzJJm0GeC8R21snU5tnX89SuBGu6NgH+cES0JOboqxAx2Vmg1jF80+1IO/jx/
iX4MMU/KGhjaQDRGe02GnK6aWan35gzHOBHwK7nWgVJ7Pz0CdzKqYlxhPCjwzXE4DMxsFN0Cr0bK
/45diDkGLAxj71YXRA4FNbg6lmJhb07VKm4/2xwlPjJKpGOs3Zs4F+0qWdWLHu7dsd8klolcen4I
60T0Ks2HsjW4KwUDsLrA7YhtIezwluYNbSuqat3ytsjVIDgX6xQdRsgB9vkh7nNfOU+DBz9H35Jw
rLZjb9tUi7buhoQ3mNPwovwrpQ7Mi0O2AHZo7NXPUKj/+2I+589xTdBmNv/0TkF2WOe6T3V6w3V7
NaanTPFlg6cSupTuG5LC19X2XoeP5SC4ukaVRrYVdx9ji7JZlXP5thLNogAR68v7Ljquuq4A36Zi
2uaIU6GrCpt6NEgdf2flSs+y+jtSYeTUk9jNfMjy34CSMsLKey3vOF6mteExqPTWpGW0gA0EMzB6
BQTUU+sX70Y4XQJPFKZHoMJ7pHMfrstoK6Hz5wUuYH5C83Vra8QS1ZLXf9hLs+PuKHgtSNAWwYw5
9A6fNJV8+j1LVLtw4C6TPIG7QDwxy9VoLpsPFooQMgaTYy7lWJCU5tbIrxY1Z3+4K2JQJIDYZWZ9
ZkYUzzSDms2773DY5KKTcocziynvWDVJxckEjofScO7Lv4K5LNv4R5tGF5uXBES5+6ijTLLUkHpM
yDNIl0usAPQSw5jApa2FItiXhANJv1yqsOOyKub8HV4osjvK84UKD7UdefFSvNRusTHl9STAtaNJ
laOJpNcphRNSrf5aL1k8GZBbk2+yc/TbV4Qzo/ii8zzAq5N9+RBwXfPp7KMCdIciF4iMnxVYHrdx
UbnvLsUd704GrecTIlyY+LbdK86ihC/TS656X8RLM2g0AzztswI6wS+gxwF25szZjDrtbXZgAWMZ
1uUtRRVwVGDFqGcu8CyNCKOlEl+mtdonRRNpnn6hAhYw2aSbAulW0U7EcpqXEA1w1NGTjouaBnco
t3dt094PlSu7PKQqvrrt3Q8fLbfD7Ak0Z2+d2tkjTbZJhybr8AhTQqkxDj1HCiMspZfOioXtl0vd
ZztXLv6P8m9arMpA/5wpeSMrcQlouV+jc1kJgzGhgMgRK2hiwezr3ccrneDQ64px7xtdf9uY/K+w
ka5VVx0o1IIVhuIVy1xPw74rVZaIrpZ4b7TpnXrm7wGIXo/9TMycNBuC0lzgltE8IQys4SDpenUq
kU6sDZ9AaDcShwDkfaX6ik+nfVf9dIToSijxbrVH0EFszYVq9FNTdecS88nHdF6JYxYwP/XL65t/
xnNv63PzZLifwXOig8pEXRMaIRjk7kimcTPrDP1yPLx9JyvleTCv3w9rWbsya3HJ6mlKLwB4vcbW
gywxtWhqGjLoQ6UqUYjKqtx+bhhUnt7ygOYVtm+miB2YQXjZpqwYPVHMuJQD+F059CQ6R/kcFC+X
Tb8osQAwb3Zjnj+ByZdI5StUt4c0//gWCA1RYuSgqVW2CRHjtr8IX7ZUj//6Xatunulz4iHr9o/s
AvXE4FgM02Zp4KgfsjntBZAf2vUEPhQZ1bQdinqMfftFlgq9/qKzEb927mySatF40roxphOJhIN8
xzxh3Mx7C9ijIc+Pc/UbP1wFKb9FHzRRPfbKYwnUvDT9sNkerSqfD88dc0d6mp1vS4QLxoUFQrZd
3FiVPoEqW+1z00DDcO/+1uam+x0fOFKJw6sj9wBy23EAAArwjqbZibrVHguYcCT6qMioY3oZrWHp
sb2FwIGPjInyskQSWO+7vlVQEadNO6J5IZkcb9KAZjL/CCFqqeFIqOS4pQ1WDRHPgpd9JhaAt2Ve
yYAYSdJefKIvwM/UnxdLxfmxwjCoWAWqvZf9WG/Sxnued2trCXt3gaIWXrfg+rxbryHnmZTh4WuG
s2C6ojdkmXu6nY3mv3RZ7hUi6fWI9b5mi5RmnmtWYplqU8acd1hQZ6bZ156hCk93MxyBkVxUEOxh
LB8GKWZDbblbBEo6OrNwRZWljr8R+/L/8IXdECF2Uv8B+PfUzFr4qGqyWPh1FmiUU/kIE0zlAhA9
oAFinPp423JMDtmzAXopPOctSu+qvYTPSMNuWvgOUyt9TGn/eyc/TAyY6Ofl2tfibEipINlXtRBV
1mRje+ZHc4bAly8AoNSXMGPZXcJLb+/en2IHbyRA8lw2JcUjklbG/ubMzVrWZoRhWfz9oj3GDD2r
xy/bbkJkUVcLh37N5gWeIFSHHR4x5iCLr+emme9PFNo2W9E+8c3A6B9OHdKZy0m2Mpb76tIw3pjl
MgDCUPipgvcEV1Nky1Wym7Ue8+3N0+MGJz094XvVu6rONksHeGGB4CghDSmR+YJUNdyKaMO5bf+A
af7yvLbfPXzPnxQhU4MUNqwCYeURtk3qYIRNkVCeNvE2Sd1W+8EyR4PzCidD06wUP+LQXSXExK/o
wDbAhAyYJHaCxJk9Ms97gbHSnq6c195RDGggD9GmrjeV+JgWwbVvK/Vlr+uNFp6K9XN7u3C5pApY
Gk1ZOFvDcRv1Kafl7D4wY2iZUOsivZiy7W56pibcqWO3peNUO//TJuMCaaCnEH45M4ECjf90GZyI
fxv74GmeDU3gfK+hrRtPYg2CVo8t2OZtMiuv9F92dq3G2N25VODiOsKCprG+3joO06N7h2BewylZ
z0n+A+fUAJvTe9zSuVSOqJG/ix1/QpcS6ICPXcRczWmFeIjEKRy3w1XyAnOE6WMRPcF3EHH3iuWB
fZ9DkzA/0wO89zKGikR0FaNd+VZdv55X2H4BBwdGWXPVKvRfquhGmWn2udx/0NjVzxxkLNXPidze
0OF9OUqWTl7pK2JgckTbAgWCQUVDozCr9/nS5l3x8tZOalZh6y3aoSH4zEXRyzBt4N9AJoyCJJcA
veUKsXSFoKfVH+fzwmZ7/FH9BKZ67g9c2TCqdEgPEY0I3Ob2SkMJ5dmsA56tnwamG07zomfI+jTy
u4dQDBnrmJnosZ4O4tXU5RaLl7sUVd/e62rbR4UaB1uqG8yH0bSk+gv3CK3oU9Xb/vFBl22JlNHH
eo8trickBFipmJcyyUqsarOtkyFALnNrZQzCBlhAVJLvp9sbuLflMVq29blo7j7xAYzofLIB53d6
90BdOOQodDmhI77vW6GWJ64U0/yLMcDNv9Q1+1KVNm7q/yRWFaoDmZdc6oIHoMS5i081diCRSt7s
5ivTqIH31w2M9Ofs6RNQFy128RVk6sd4dnTm8zCfsCnew/BGDP1QOrs9IC6XBqR5WTtPcnjM+KJt
E87RRGsbbANxbCBAaEd+CRnxMznLMCn3Rh7X0YZG4XrIVfCyUlfjuvLGJ5+qvu1OIHF+TLH+f8rQ
BpTEcErFlGDfXFDcU0FfISZ80FbcDbZLMpmJOct8sCjl2/5iIrRO2iJwxENE5nHvtTdXN3+KCLwh
Cnwtbt4f/Qh0Msuiy0Lpk+2sM/YMtnoXZ6mbIKvz4aYA4wki6AHxCgpuIs4qJiyB/8YNEuwjBpOb
rmPUSWp9BEYnitycYl3k0T4OeYuPj2/BVvNRTsTdY+m3MtR3ylSgatFEakVpbg5zVtAv2b4f2wFo
rGCiPBoMIgb5lvETfPBD/kfAIw0CWpFaKPAwG3fLK+bDGlt8BWZYUeOPZa0xMpVMS7IKzxXRsRHF
//PZqjEILzwUXP4j76z8AC89Upw2SWm4sp+ufLiIOLGU7OuZHWA9vGlCToBUj2tBFJ7Bivyj8H13
QBorCnhL0vTeMHun2VDtCn9Q+YELQ24HCnGPWeLbZvj5WCfB2P9Xy5VbAI7+8dbw5u6cJZEWum2p
UHaxOqcEWOHK/GuoOMsB+34O/gDKWf/aFyo+QqVNzgXz2f15IcQiLURtkm/XbEuirrLFj1gmXvt6
0sZN/Ujg091G2hr/YqVJT0orf2ATPwTbv0enJloYHgotLsbXkxJCYyHyFJhHuVznUSrtU/NL8PX7
kAZlRA1ZjKMJrR22ZujD0Mmlj6ymqHpfrfOxBKl+7nHLcWCnrA3mdbE4ieXVybCoKU/fB+8/J06T
SGtM2QLjkkbJ9CsEP9PE2QvwE3ofHP+gVAz565P1CLlfZhpEOftyyT8V27yRF/uDy00qGqhlC/ye
YAEfWzc5SeFeNPGBPkyXw/5wZ/bgoPrYgeY5hKDPgQZbj7/v/CyYdDUfmeEDEhqwfQRkKypQUTz6
caupRbaXAGBBnd6otK8ql9cKFIyzckXA2H7INSB8W+0bAKEfhnrFmvBGdguuvh5DKSxH8pfcHyHU
gvQWqlaYobiDh9uNUeEQcyMgBlgiur8C4jwFPsAKWnYMQsAupIdACP67+zuo3DWvsl00tPqRcdIn
Vx91bNLZo7d1eNQCt4Uvu9Tt5b5Q7If6oNcx1aG8Hh/swcdX1986qmcYya3REYYVzFqFfyhFsIj1
3TzooQinX/qvcsgB1wGDfLcBiUL1HYmHtJEDc4hftmnnyVsvojJaAeBGh0xxPpj1rSCuj9umy9QC
YWCsj0BQlLxl9RrEoFO/lzXg0I07R29ZadPw0Q6gmWhYnG9i3C3vKPxO2eSTpB0/SuhSOmBqIrE2
2Sz6l0wHHC4140zWtRuGAvGjklUaNnkFEiRdegrcsRmU7JEEOIjydWDFq2VvWZmcr+YiSlnjoROD
9ggziNTxjH2zePEs/5RvpU0jRdodn01W4ls5+zDMXPrOxkq4rlt6ZZrF1Bgbp0KqqLQEep3tVtds
aQEqtEa8/geCLvP0atfcirKpiIA0C/Q7XahLlMswp32kgc1Hm6w6OiJ2fXR1I3SqJwd3cicIRv9j
tCxCbsuCsyBiy5L6mPfo8QJB5SeKVnMCz8lH4yQJd6VDVAUppccQ+ZURRXS+KSicWmP5LhTIToqJ
ubjwqMhUj7AelAhWAAFll02s2unUOZEqgip5pLHtxEvBdgYWJ7C5QlRSYEllE8ByiUPFGj2L6/0h
n3LAOS/zxpUnmISrdrRIqP51ryQSOgbDDpueRDmLheNROhA0KtUBvT1mQte5D0MfnjXoOy0v43m7
uz+L0KhDj5wB1AV+fH+5FfbKD4rrJZjsaSSZLh+SnKppx3Y5JSypN8ILpnmLqU1YpR3ZqlxqeZ/J
9ktfwdxPXEDEeorSMyVQiLw17wWyBkjspV987FfIunBP0Zgm9oUIcRWeIo+vBBCPF4JpR/oJ1VhA
g8vC+ljWzkg6AM1hwfOPKvz/9Ob/wheIlBFhuq5CceMeKJX5Ip/LtlXOsOexO8L6/RvFklCkpZwR
LmlFzlBV6GFCnqaGni8+AxcD4uftThn4zaMS+Qsd4or1hHHv2y8ak1m+LNKDzFs2rei6O+FjmLc0
/A8hDhMUnn5pGZX+hb8c2r/sqQjNZWLvZylqgQ20mWZVs76URrxlQ+1glqjbxZORUe50nmG+9M9y
IW3qKAWe+Y4DlMmbeojGv5sMuSPn3NQrCcHnJP+7U08UJuRcIz052KRjx1+1u1w05u35FTjCLtCl
BMomx8RoJsrViixa1zw2h070CX+0N8H+n1R+Z6ekV79NH5e3VOsXOtuqaY/5mWlljo+OOVhraaGn
bvjDVaBARHNHN9vl3qdm01TomiJCGUPsSFTCyE/vvSdp0zTgVqi52sa+TsLs6sE1f/2J03aag8l/
NSvroUo8MutyTVTjWDHnBgVLXslQxymgHrdvUOrpLo1JKYowAlkLws3QnOM/XX/Z5N9Jm9ggVeZy
LeJV9plwtGhZNTBAu5BLN8OCKeeX/rcpSK7O6aSxW15x7sCKiQrLeaq88OKWaDHvxJZUMxZaHEEj
Xhzndv8ssCVlTHR+US9JcwWg38FOhycW8Iz0d/D/41dz0ROWIntjan3sRdzElfNSm33jgAnSL8NW
TU5QMU3+FpgEsfDBG76sJSDNRJ77oB/O84E24EX3Y2fzd1cQbNlZz3m78VlQCVcfGnoFzBnth4JK
bOAR36oBp2S3yFJxbka9cp3FSVODiUIDVfP9Ya0Ez/Rbj0GevgA00AVRJYEilvQYQnqSGA8JJ9yF
2d2Wnar1pbtOuqkYIflr8Nl3AieY0luztJUhXjUySOdSMHAgPelwrlvbph/TVYGZUxoqIbJsUtlo
lmrEESrhYj9fo2J+WFJo+nFqQ59mPtJ8ec5RIgZts8uOhwWgVv+5Cpod3NOxTc7tn1B8XkmblXyp
pgIAHa9iOjKFKILi9bUa5iV4GXDuWaXf1SIn7hSxL7OsEdA8k9GM4lFbQs/F94Ltr1QE+3Zl/vOn
3UTfj2fHjnxf8LT+NHXlsYFfaxVzeODo+qcpvPW+i/RwOJPbbiubM/Sr7cEOY8eeRjiIiMGkzlzY
wTvFNz/aoqe8D3/An/RDfMpZMvPhwWWQG7Jks88r00qNrJwWvPzw4YjKCuMFWXdhtrFwbfq+H4ua
CMKCjzqFv7+4PT/nt5XQyEYU9cHWdg/YpPYroxbhFccbW+9PS1cp9E7peSB0YBfxJGp8ogjkgkQW
YITQ2MRv/4HdNRzk4FWhj+lAWgTHDKplaZIr6ZTawVW/TAr00nqIuo2rvyUxtqLBqPASw4eLkUA3
xKSTlBNOO08VEn0RM0Oz2NK1+13wKXZwlwXNFEEg9tKN3LCPF9om+brf4sjaQJdJonmhYqOqV05l
VCQ2NocVxW8KzDEQE9j2mkLlxll6ukNd7Ch4P7mOd9fX7hsBUZWM1WkpaE5QJoNeoUjbGacnH3se
BmsZtEUrKh96taQ/AcxYhpZ3D2viJFktw52Tcpt3sBFf8b26nu1Ngu7g13yG82jiRUblrf0Nfz14
b2QI/hEpmzxMoax+/hhj5ACcd718ZpDfy2foAkXAV/JROzUu8kH2zOs4kdsWrShNso0/GEvzK0zM
rdeTdKcQU4o2OA1dmDUYPQlW1gS45xow4xJ2svd0990oEiTbaQKSFSJtHaucBgvEKfGB0fJbx7Pf
BUUGWHHTUlvfDpr+PW5cu5Nv9c6dCFAyl7aJ+/n2dVTcVnFloVVKKFqYsR+A+cKRVNblmoBc7Yf+
Au33X3iIxQR0KFisxDf4SV8paGZbf49VTFp3EaWQth60GRXV/kr/+MgiEAWrzuhfgeIQ/fghmxIb
XAqK+3lqMJho+Hng3ixmkqPVDk10KFnKQ93AbY11Fx+NFVs1CsZInH5oRUDFZfnUFRcqsFtO9dA0
nKoHSQA71GDRh1f6jsF6C2rV4fNEVXrCEil1khtjlzc9UbupAGWz0pk4tfngI0UxfZJCqllZuufC
8IiLeG8pCW7QIznReL5R4gBbAE30mp3AITH+BNK3tD6iSj1gy+DFUOM+xMUXyIMwkXgXfoj8vMfk
eCvuuWqFqtX5OXPuZdj0FXZgg4KqmA0xVTjJZzx3XPFEC1yK3sPOaWdAa5ZRkXO8qwpaCpbezyeT
xoVTjUoKt9Q3xZTLfBnO3y7dR4MSw9/PbwnbZxViFMJyU9IS3W7vJjNx+t2jL1sdKeNDZNoMKRzC
9XbfpINFCx7UkagaK75sHX9Y6GajYg4Y8ty3yF8FZ/FSNEBTFO38bNzSKalS+H9fmfMFdS5gezBG
4Lk+Nn+crI71qtNFyGVHyb3WuGYFbElO0hhaq9XtqMnyrmarqBc4Ez6tlH+F5Gs6N4mkHkqCFmQn
BFS827OsOttmsE4HTL6/0aBKqA5uJnSHY/35y1YW9fa9zgH00N5bL9utVPGnqyeLAdJJLaPOUOll
TyiCWwysGT5S2RuLMsUXANYLTgF/qPgbSQT5+uQVYNE48KVF0JrIyAPLRtyVTYNBUahj9YMhgIWc
hUlh9lr4m85xUJiG2vX1f/b9mheBw8g/N9aKBdvXCDoilbjAP+/kE4dG+NYo3l/7LEIHL17iEUnc
UiDKuek1dn6QRLTG1XLrzAKaL5tuzIweSsQsI1jpOzspJd2D2SoL/71JDbi30fwtscRsjXliW+st
gXHejM6Oy9AC94vVbfZDo+AuG2pBAWmOLu213YJTrF0LBs3cWEM+um5ej5cJ2wRoEgcY2By1i2Yk
DNQXaOmEKS/QzVMcyTqn7uH6rsIzq+yxezbg4W2Hr+BvRwC0QDqyQ0VH8NCQJGbBbMR4YyVwoI1Y
cypMksE/OfmwCwej4Go7MWJsa2Pz5/YvGgGqPE1qbl9AaOQ/hSgHlztMwy7/WJIHLtkFoGSoZNJb
BCLLGUzPkYINeKLI/ofz4tTYF9RvVM8/MXMolFCtSfdfsytGZ7yPGS7MisN7v1X0tB/SYaK9MjPh
M7t91OQLFXNVw5dQs+c96GRULsLFobg0CIahxLk1RNoJyhjWOFC3KIUXBnRyI/k9KWrVlq+6/Y/+
XofKF5b1ffxdOd+KDywhtHp7c60/f3duIWCi0DTJ6sU/8y2gdkAyhokcIWfiu9aG/RekXKEfo+8B
i53dOO9ftZadWTVOXhuaO240PrYGr4Gs+ERdUgUNkJA9OJtEyP045uafw7OL0uoItu/0lBZLvcTl
wf3eDoCSy8iENugWSJY2bqJBBZRnQBccXR6nbg+BLOixydhbnPRj79p77ISVSNu6mCN8vVh0dI3c
/3iMPX7JiCnG+cyEeFuvYNPpylLWyKWnvQRm3y7QUaYwnD1cGcFIp55S47qm4guGTWewaCo2/TkI
88cVFl5OjUAsbczrLvSefcZuHYSlv51ydp4wP6bzaafMMIrGBg4AUDj5iNQJLDy+/eV4OuoQyBC6
co3Ew+noAi9AnliWlSPsOfnZX+fHiKYlPeDg0qS365XdIQ/beR6TFdChsbnuSYkpa6dUBoZNg1zV
La9A3pjOP+AC7sUPDuyxiKJeHD3lebzfcv9FGulp5uDEDsiHpzyU+N6EQDW5XQdGcpXy5py21SdF
M1ax8S1ksgnfYtUNY97CfF3bZCRhf31Vxp7yWdyMkcr9Zw58r2fcflPcKH3+IyIYnSLNm8u5ISRx
6WlJeo9x3D97DEKzB/JTBpH22sY9rrIM20oSfnIaXR3KwqFd4LDozTipFQixbY3OugTe8ZBhUbtx
Z8qeFfPNt3ofiGJgqg9GRNVR3lmbGV9M0He5wfc/mXzqkEp13UuYobMDwv0jWVfXC2C8MJjw9/Pc
i9Eokw9RZNM2NkbN0S4RMt2UpsyATzyoXcxS4OkdZJXlncD5OOBYGLTbInA5LHp6JxGy+WqiaM/h
/U6urmIKxHilSKzNLpKBN+b/+u0d/EctxMdRDhz85a4dFmzdash+QRzsfdA1pjl+vbFyTXTFrQRP
EME0mePFTslYI8BQgYK1nHfCc/Exwjrn+Owv0QYj4miXwJ4TDd5oPe3uBZ7tdnUSScI5AjvU/kxW
H/Hmta3sURysAckwEptS/S2U7m0iu9k3BNSjUutsYxW72XFFjX5zay2gg7RJIOYR+30nRIXi9u+t
QIoLEdkfXS0a/0eVTV8YsPsDoufmR39tMAhB7DthtjYcQFrdC9TNhHpI10jyAa5luFqHyWuyon6x
2UN5Q8SMESMvmDIGiUFVVO5+bcM+FZlAZrw2gPBCmEOfbyfVKfjbnP/J7uyuKTWCKqg09Qz3yPT4
5+aafQpXUZ79xVkddp0MTQZcJiC5oZJ934w7h7PN2La2J346IwRV8AQi2ee/kwNO2UvRSRUps5Uv
b+GQQ+J06HEKxPal4gKVdzujv2D3dYqk18Hf6tik2dsblL8Q20MPH+MrzcAdfBRZn+zdTgHsuezk
IRvzgQKle58q94RSBRAtGUaXq1rgDe32F3Y/8lxKCWG7FRS71+0jb2FqRod7i33wJDpg0yACkLdc
+w/aPBu6vGkgzWb5VygGu9F2C557Cry5+xawo3dv2v7e8M8/YiEiebTC7x5vCzvH0Blsnm2Up3fl
42mYr9G4KJQNtSPnds36RjjtLZqrqa3GOQU58TADAFDbAgj+bQRsb8Bsyyg+ZkJt5c2vdxMg8cYV
uKz3IIqNHlnhDxGk/ewdwl9ZUq3Z9Cb/yLqeL9O7tiuIiW67XF9uyPgapJ7xQiH7WOK5yReI+9vV
PM5dnKbXleVEs04nN4l/P/tno7l8fl2ZsDZ/woaK8Aa64jgQMKyUg8bz3HxIVxhyQzD7oCoZgRNW
AFVyftDxXlAOX+qMDGHRa5Q5pBMvOSdL6UQc2qOu+2oiKxOoRXETywHnsqcB84PZhNs84vt4pxjF
j7MyRyncIrSERyxEVAf87Ae4uV1oUy5keRZEtP6/I5MJzot/Cek9xZ8xkp4EzsOYsawgKf77mhWQ
/Ync8oTCDB6lYhXaHuRAMRG0VzE6L7/lBmYcqCqUCRaUgN7F6ZL7edrVOklPkv0vdlZQMXudwhcT
LHEtBXB2wMXODy2kT5pnfJ0dHpSh47cfP/iCTW7DZ+3SDNc7SKPbKaD1rak6KBvtvJn10gHedHAp
H7ZTpyANC1kHTVeOupBIHd2AAHeC4erezCNiuPWo5frzWMudiJOcaISk+Jx72+AiT5hrXj6KYvz1
qqdplsG33NfI0LSOn56B1jbO0KQJTlFLoWaO6C7Vo/gFb/j0plrbOk8JshjKNkie/K75vMhM/v8M
MShfNoYTdNgTcvUxQjHSMSuYgEnW6+CU02l7xJrztrGS/eFl4Fz+TS7xnPqf/V4R3rISpaNQxOVy
SOrnyATuaG+wbg8HVAenl/Gt+Zu/JI2Wxi7GwfUnkXg+rvxswPd+bWVQ5K/VR5Zh0TOyFL8s0pkr
Jtee/TxKYbz6CwWzj66yTlzDyJEl3g3MmnWDyO3B6vnGn61VUcFF/XZI2OhY2S2fbWrM8WGFDbiT
q2xwWonMluiTW5P+cw1IokJ8P0zB2IoBqzeBpS+OJUrTZy6yjF/3lYIjlQYGGM8YDxnxeosc0jT/
L2xTQRpd+efYWVpwqKtQ6wduh02BV45Fvr7gaT52Rm1Da6ONMcMMsJ2kzhl1cvRUUfNXrM6/1AEl
TKyva4Ps95uddAus2YWwXWzFEnHTxfP/CTlS9FzZhIrdPUGVdNkcgrvM8r4zB28XZax+CrpV2uoX
V2OppvuNegikUCFSA42fWdAINZQzF0bnf7ihLpgdYfJngR//ZCjlKYYSiNTsOgQIKPi4cmWhkEx4
iwko/0lSiXNI6Xkcax9fxO0kmIWImn9LzzZ9lCaSj0ZmmeuWz6PGCAWR0x0RhWtCleY9uh27Z8pu
c2euH3mfG66jSqIzapbwJ3Qte5J3cPk/zi79EktE1pfFRK1cFRtc6woq3f2JdHwJ90unMjYMgjmQ
YVJlohWtkT2o9WEaS8f/Ic2FO6eM32tcA+BSS3n92aZLR5rgfMTjkavT2d0Y94W4rkHnbBzTKG/8
3AAKp4jh2DZRsmBrHtIGHu+z7kCgITeU/d+o8JqaE4+Q1gN07EKvLWyXfZsBxPOQfdOj4xklOifD
kb+BnszVJSOXdhgrZYCo2jVfdRl6Om+u31rJiewLmNa8XZtRejBtkY0zLcrCXHEc99W0n+1yneDd
f8IT1Dws7qPQfQxotJ0JjK+/yqGRt6QDS8cs9+zbOo5aro9h4L+T7P1fzY3z2EVe8uz63ClGrFA+
l1pk+EdazaoVyd2Y7p1iYfYVpPq2i8DWzAXxGOIjA+vuP1oBwkvmnoF1SJriN6dDaKCdgEYwMlai
0H/moUVECTzTmRXXelDekD3fzaOSyEzY8pLiNQVS5D1TPuYKQtrK3p4K3yHD+CaavudM75A/Wz0M
Qbx+Uf9XTP63i/vTMjFHzqHOy0kTErN3Fy+OpI802GxHl/VopM+j1lxW4Nlsy5RKKzdVMBGH5aOF
HGdYxlBRMpd1+y2NBO9yAtLjtRi9sRdEI56H3qkkhf2WYCpCrLJ8WK3Z4rvzxtWJY+C6Fo8Y9P9l
a8gl06a+oBJny4VVyHlZd9nl2hIaBxhgLGW2Qj3XKlBfffB2vOsvEtYAQPec7wwHJYiXVLrXjweu
oAndB11qb7ueJoUw4aDQXrBwqcQzG0RzgLTpvwhJkE1L/L1vFOfJTM3l2B8OVy9KetpvS7BKz3MM
mSsOBr0166MStuE0UE8ofcszWZr6iUFWr/52BZfMWhmKFC+PPLDbVfNvBP3BKqpKwC3TgAK2Nehz
S/unloUycMC60fQsh1mrg4dsx4O1qHowe8eIq9cfLI27bbZxEdko9lWyjHjIXCkDt+U10mc7WgtS
XybOd+7VVay7xOWhUhWRj7hcyblbOTBF4dvcPEtgM3Z5qDJmX9prg6x3S9TrQF8asp2YRP8qcwvz
HwKHXhPAnYFtm/wMeSykJhbrs7NZtD3Dr1p3aNs5dGmAq0Nak6nPlcQ8lX4RZjol/pGpIlJbmHfk
tQQtgQSF4+VzxA26LfgZS6rs2xrlNbe4qjBnl95rrPWq/tOAeh0fa7eSSRBFeLChbl8eFb1U5jGN
WhRv3aPCmhOZAnTwGHaZfvZoMvX89xdpKwaNQ0OL/LdOsLMZmiASMa8n4JqagEvtqkaIJFF44EqI
Z7BdDD9xRqBsrcJgeFIjKm+gKnNA/oGAYU43NSjLpDo8/HqtvaPy/HFN2CqUQromzTOzvZFQq0ac
7NCzlUyeJrLSKj28xlCBslSLLULnsADRa2eWCEUXJ713SgolNkQ6Yi3WdzNsUbreTHOzPuVN/1WK
SX/Kyd+IwYq8myY8NfL29RmRNN4DO7Gz523uxggIlXqovhXzbKoahMvtU+ijG8yr+QUkwwL/cb4c
XquUgkRKn8RVFfkAGDv5tqBtDkXUzXUOqwIXRVonmOQKNV5Z1vUyPIM9mIFFcxt52LRabX5Kq1hN
uihM/wCORHb0Iejpx1MLAnCyuAS/ZtF7WOGNF8JGmx4cAUj42cXfzU13hDeexAN4usUP1b35+vPW
E14mizGyifuvC6+oXO/kv/pnLXk6IVqnIQEQkt9vwgjdNiEs704lsAjrSGIP4LM5kCIx3E0wtEud
onFEN3cvBr60RR+mOYFDZbQABKiB8HH16ZG6VrrWDAp53nMBIxDvCbTK+t+USjHU2UgoJThQMxbA
LNrWItfPGZKjP2aWyYIPh9Vr7viCU4P9tEN5uANIp/Y9ASV50l/N9/T2a0RkUtLiTD3tAsWUtFOz
vI9aB41Bdhn9IZvJEP3X8g/GLKqwDdClQMqV5g6GnBqywt8mt37b9Z9JkvPpDPbhkyLtBWpVUkfk
JRWt50yct08KNm943Fxl/UunUY8IuQs3063qNYC4hRAxxUCF6Eru4Dr87lP2yD3Z9B/toYajMg8K
07LVPBdHlJ8ZHLxIo6Rrmt5aXAx7aSCsbfqPqq5d/ypTRG/rKVpCK3fAlFxcVJWcfOgxEysYcH5Z
zC7TmginlChtb7GzZmwDelc1Piz79ef3Ni2yASntFi48EgJRNm/eo5QDcLSeNFVSGhYcuRZZjx0A
c56JEdKYKFmdBqaMHCOeatvdL+hKkcancdPqOZpwszYJcfEPoyQkMW+3N8GmeHzVjZUCsINMHgn3
ixGJVD84232vn9uLX9fLbw/w1cLLI0wYQPgHLfsoJReLty1A9zEEpX7j4KNlXDFRWsGtU/aoMQvY
Uj9QJQ1zAQwIgku0vanIV50TL6+//hamwS5hIIhx3go/492UaOmSzMKHoj9jETGIiFH1k74KwoyF
7D8I2xiBVL5mZpGmTLvSvmGjs0tnI1aTp+c2QOWdJqPsqoW0/VHtH/K+8/BS3CewqoLKKCOnWPxZ
uVuq6X9fDJ0axyXpl/o8a33gAj679z+wYtNoTS885iZ5jsdeW+UruoL7vYnKOn6aq5ufzuhig7Nq
2PlqumJEV1jC5X9hDpwPuc9XgXtk+RDJ/LesnAtYANP3YLvAazDmY8XuTcnyRGfYS9CUNREz93Da
5ykLaBcEvwh9doTN8+dUdxZwNBDPPSXiCLCdNTwhdffd5MnJKN23wqPA6aPeVj7R06JIkn14+H1+
G+UBD3PVUltS8KMEl+TBKfKKFMcCssoPdkHII0qTFp7RuZukTi5TY+cxOxrrFPxDltmhQdS5Mbau
xSgEy6MM6+MLEaoKtqFe7mD1QyJiUc08tcAanhErxCOhI5/CWSftH3cH8TffZdp1sX5QbiJggLHq
lJqQnXq26XjXtYbebQtL24Afg12Qwc0er3cv4etYyjxQ/glX/p3EbdtuFoED4RvfC3n4+GXEafaX
noOPVoAcq39eYwoyHvtAxvr7/qWQ8HIFXcvPAQTBlYJbz5+K2pwu60rmsKVD0i8NU5mQgIGFahpQ
evlbZjaDSOpWXNstPXkfaRwe+Fju8Hk1/Wxm9eTpZVQQYvbH4MVD0aSV0d1E4zmK/BCgyZu4NJAT
LQry+HmLSzSwrnY+pBnb/yjFwYh5FmyvKPNSZkU4O9oK5cKcsCiRxSLwOMs+iCKQMFRV0nxJ6cX0
HCzpl4/RstMtUSot3E8H3W/mxvL4vJ+ERPtfAcdjMbl5cw+Pb6OA4yEEOY7byfxslXmLBFQa5h1Q
PiOnSI872zoTedtC2c5r4Np7iYoaM1r9sGN+yftMapekn0+IQ6vfOxoicHRMvTueQmmwi8Wg08kE
Ap+nfaZrrUC3LtkY2hsNQKG3lQG+kOWfnQuzw65nZIgbwyp2zUdaIQUsLm6Db0UhOKKpu1bFlp6E
EHHh5nPQa9F0K4emqXpNTjAroGAk1O91V0d+x6KDZhaA7f47y29TBG18CLUqwChScN4SI2U54ZYj
UKU/+xy2FfsYcxR/yvui1eJ3jhYsg2opr2Au1a8Kaomv++iGbwml+lBElCztOXnH7a08bX/4yXFm
/L22IVA34qf94hdj/j5BHQTb8i3Orp3AXpX7FawSEkRXoX22IAl02c+q5SF+5AABxb3eBvUdvQS0
J620kdM8ura0/HVMa1XasNjtf3JsQF8I7WIPo7T8aTvG8jFfVzgc1zXB50roqVS9sYQgoibdDyH1
zGj6hmjM5WABwTol5nnpAVcZhO7VptGuXvrZOXcKyTD6Gt9TPzuKukwZAqAsgadtJTn8Sk+TYVCx
UZY6PBsYVyMC3hQ6jNYgX4SvzGCjTf6JURoSRlGBzcE8Du3bNO4uS5ACGP90ymkMcdY0FczORksN
yXx9NxM0oYZLjPVt9PdmRUNssW7uito1e56SYms4GuIO2D/eManMV8uY8QcYhp2kim1htiGsTz+r
mqos9rIlg8Qj3T8HdHBlhskXyB0IIScZ7WyzRGYTlKWaMe55KZiXSdw47ynRDyx9jl+F7qw1WftZ
8xTNDr0F8djUHPWAYAuNFK7BMpbbnp7wEH/ANf338PmbcBL1VWc2ptUMjE4o9fhZyokJ3B7Y6Px0
M2NT20YjqJOeWKbdjLsSG85fx2vAhJTwmkVjGiNOdrmvq1YdH5KiuhHm/3wNRr2ADdL74ohyUaAQ
6puMWiE9DJfBZUQ6o1sdijnowMSumhDboxdywoEQMaicoVRd8lvSYR4IrRhu0BDPt5F5ETvpWpOs
BCvJAvqF6ETZYNyz41BkqSfSrs1zt2q0oyzB0q699z7cuw3SgQdtUEz1iTXDYpDj1OFvu7b5+EdB
MBspmKfundwZISQ+jBd1eSqE5UduyGudp9vIb7SVVI2SXTjGoTJwQ6euhuBtbRJQMD6JEyLi7sOf
rTpx1OLQBXIPzoavFf8Aj+KQXmGU6rfdf2ydpGe0aksuEPr3na5FtSDjeZmlc8k+4FpP5MoOcjxh
g6kBziyjn4fRu2SW1sKld6Kf0AAIt8IF5Eu3srGtERGxEVUBb06Um8NsCbaxZi5ZuGMvI/ggvxe5
cqgjLNWsj+Rf4Hj2OUeP1aDMy/Uu+6sY2JsReczTApEqaBF2hjoJLGULvqcwjl1rNxGxgaImWG+V
+7lS9wX5I1PCTzmwqnjEFATyJ1wgPKhclKJHIlLcJ/pdZfHeKqeLt0fPu+rAyKasMpkmzxT8iOFq
D6hSUmlxedVxfnxKwuo/lHW0HcMhPm5ouioZRg8SkDmegQCyU25wvrm0U/L4AoFxGqbd+t3yvK9m
R93OBWTeupnYewoG8o106c+KcAzO1wUZzha05oU2jWfL6hQhkwpxWxpBTDD6dJS9mfZ7/WpOFRxy
ISB8NUfxKdRIVOkVsmuFAw7LA8JKbuq3z4tEjUhg92YoeCLHnXn3v/ljswfwCh0NAGLm5sdoqDOZ
zYnZ5XpZHszNKuHR1iTdkky43HjXT9L0LEJRWeLL6Nj2JjAZhh87NtItg83Q66RwFaMm9vHnLvih
eag4qSFViQpieVt9njGTz41TMAvpJTWb1B1P+mAGSLCkLfbIUTbEPc/YZFxOealP4tQrqdb6Is7Z
JkROJS8OU0WDk3FYPvVqa4WxtFMvcOm3dYyLDN+8Rqi1BOOzzLzEPwD1s5XJ3ri5Ut3Gdnshm/co
4wdcQkK4bbAp62j4Gw65M27UBsqKG4ned5/PmogjhaNjbZHHXBfujeLjo77y67By9/JTqiSsLY97
jzeIsYzkCpJHT6ll6FIe5tU5ekaA07gMUCxKQIm07H/bJWGO+1wGPdyuSShFmHD6hJHPGCPrR3Iz
F09iw35SmljUkoRtqzosTa0iZ5D1MTkJgu2rJCNHGaixKWg+iXU0IQpffbydgkCnLkBqk3KLFKNh
nnAGzS/RV3i+ErIb/MWbRpWjuW7zaB4Id3+gtGZTfGFmq16omMZq94bAyUHA8cpPdS6WzhqFXBLt
m57MypmRC5HIqhfKlaGTlKuYhdPYr5NYMUjeUuVbKt2zYIR0BNS/YjFg3MepzxNDqWbqFqVBSQXc
vF6GtthnBX4DrILtwhMuVgypezQd4jj36T280NPk2LjkujMh0xsLyf6p3LLB6xnIiBuqpWTHCkHl
PqU16edOGUE6ccG7I1ndaO2UdjWjEs8ldhumxNBX0YBqy+gqqxWEpbGqc7y4+uORZm62iGVhGzTt
zqrsmDhQuXXnijy7jKHWlwaN6oOdv3cMh5b6wpmgIN3cpLowJ97649Ob0X3gWFJYHFioDX5EAm7B
jp0jBXBEJoxN4bx7VvU3m8nEcdfilc1pzoQ/44efN4KgNvJil0khg5+bWSnwsqGZuPcrS/X8AcI9
REQhC8Txf0qjOaFF179qladLtidMn1+beNOZNfP3l/pyGm4oPzglNOKvfLBqVxUOQAZ91JT/HoO+
GWb4X+cHqDTMLSexEl+xZ1tcopF2G36hL5LmUgB0kyL60uazTERoUr/60mP8bxQeq3IZpF/QNXQ2
n1MC6JSf07ZnVoNK+NETMecuuhj/W/rHtvq0lVhLi4uAZRLuSaKRYDtbi3ssNBz19UcshNRCCLit
k4DoY6uMrTvNfqriEsKA9WzWZEU+xWROaUccczaKsbGvqekRf+wLIUL0M3IOtEIf3bgagxAajxT1
nHjWmiWLc/jzD/EpCwjhpb3pbFsdlsChpnMp2b2byUTEOJEINk9IRUkEQglmzCL/F0xkDloMD0l5
RsNVtxCxSLwqajV7zjPofYT2b4810KSADo/0WzebtUozLILo7vFXXCCT/FJ8Z6IIxxQpZO+z6/u1
hMR+VelA4ET9OnmmzMd3XGhGahW57agrCWsAiSVkzPNJb5eIerzvhhB2unCToJHUuHyaAeHEq5OP
yQSFciqo6BpXWzHvZPxa/8HASlrrJqDuc0FHtQBti1Fn2gGfkfhXIjSh50S8ip0erOtJLoAFvqNf
ImsyGA/xpEqvk/muAQLGJPP3qyRoFJ6JMpQ860axyncoX39FNyoitDacGxYe1+G4PaBR1/kEJ0hL
iI6c0CQZCJipNAGqRFHHKwGKfpRIkOjenjQOd5rsiXfXcofpymK23xHyAtYprcyHVEHk3DzOpSrk
dKVQrijbSddYDeNMlNfCcTUTt4bVHkwEEKo0Kko4us+eHQzOsx9Q6VTbLNE0VVb4A9sEOcweeeKh
sIYrbuTXGXDA0pAlTS7dsbn1HnYVYLtvsbzsDMkIo2zc50RRqo8uaT7TenjDYKiewPsOj0y2W5Qp
em5eOiN6GwKJc9Ybc+wxfL0dg65ahvOnvgGh/kihcEFGI6WPWqPKd3rTuenjZzL2CSLtqAzlxroR
fdpLDnfbzE/GPt26QE6/Lr9XSq1hYaiiCvcl2x6h9qMF1WrStSQA24rWNBb1AFkobYFPYrWBCEi7
rKDnSVIphGs/HF8Pg3Xm2VMF51rrNjJMhWhz1PMeU2XIHDSYaGXO/S387sdstuCKSoUHNtuuvX79
6eaJwqhd3wyM3d9Np8rZCd/nxAXdpcBQ11ydLnkjRtTkDqsXKOf+pOqacgzrNp6m8YiTgpFEDqPf
LjcUSJ9+SnPKsKLei8HNya+A7UQUB0FeiNkefiZSweiZ7Xj/ODWNPJ2K4PiM/JtTYofhGfKIzw6p
DkU7w7Z8NspSAadqyH3p8Xz60W/Ry+jGJ6kMDtUsW3IJkHXs3lKwaKhteS9oOU49RG7lONQeZ7UT
YnWvgLOrkq6uYUmnneEKoJNeNOb+3vZ0W74joDMbe0cqRqhEsaV8TBCQubgeo3a8RjNa1jHPzaCP
yPGXBj7ofiEEy4zmh5s/AM7A63Vdl7IVzHscOqx6u1TXgWfZsdJXTpQKS4Mtnv7HBC+qeAsiRd9o
7ftEQ4AcJbRq8hqqCpeXdAs0VHa1UV8i3FVoRvUEeUhMPTLF+bJ5CwuJzfX3FjH5XkVMnxkISmko
RFR1+FjqQ1pi+73nsTVT2XS4wMGqJuaHZOJ0CQ6nJuR59JebDTt4oE/Qq8SK0QdeKpU/NlAXj2es
fEUpC5SYQVk3S8uuZ//vzWaaE37D94nw111Di44tWFdqY2gFhNkWOt/5ZWswYNVvE3w9Lstqh7Kx
OOFMg+FiZCZARNOfW+M+SKWHmkRezZqUPpV5D9J4Yliz5LEgSoWSC3HRiPB4aHUct3xlxMJLiK2J
gN+nPuIVZNwEWpnV1xf1ZEsH355f6qjq+2gOZbQXkM0XWXW6lQMW7Mzq50tqZZ+KO2MqMI1LopOb
wwHYXoS4e33y236kcWwwwCSpSEdKa9K9dmvkG5uBS5vjx7telTp6KEkfipFFPJY2Gb4IJLLZzr9P
D1CklJ139BFFuXAXqVIH/zc9PhZXbGOR6NWFOtALx0vnIggx8FFEUjD8hedO46zon7EjMQzrfCdr
1yoGh+t4RDsOq1mCLGC7bG3ay9lICDGs33VzdTpDA+qA4XkXBVlqIZ4fVNwgPMQQUEu9voVO2Zjw
+Rn3T0+YH4c/l+fRzS/Xxv+WbGOAanbSvA402S/3fZaA+Zq70HiB3RKFkrbpzrEpwpgDuhIuX5jH
7xguP8cGrwluBc7KqQizoKiukpWitl4qyxBfFDg97Cx0KXUG08iOEAhg7o5UJFsMXr8aSHUOexX4
XPSTQQ004qZyOEjlK50ABM0vTl2ydSUYRKn2HGwFzgmaiNxXuLBlWH4uexcBIkdR5/Wobb5c18HO
mq3nFJRzbVLmJjlxd8u6IiiwbGPM+nZCci9LmwiH+Fa8Zdv6005xV9xrBGGOJCoygwMNKHCM7sWc
aFDi5h72nVRB5H35lE6be+iO9CP1a477BL4mBpHvBplZ2uvTj8Xccf2WuWnG2AfXfu/YNvPNd1hC
K6TmIQ9jv1lLRghndrtsnxeG82Bd5drQ2p3QvZDd+LBad81I6/O8tV4+ZwdtYFVL7q3B/qtOlV4J
suJjrgRF19yldF18S2UWlW4TZgy10bkkGXpU/uXOfAH6Nf7NveYUCBqKnOp8YqZvaD0P1vhAz/L+
3w80fSxUIKBnXEksKva0eHnJeVZPUvu4D6J6U0ucUcDiCFgNs+zDOWkh5zQILgyWwJ2079w94XIe
q8gwZ4zuX0A7KVW3uGSNBbxPFGZ8mXD145zbxLf5ogBUTeLjbRZYI94MfNOdR4H9kx80rzuUSMQ/
eBqe/abNXM+vadRUXzh95uiOEtYGqMeLdCXQTc+cNpug0lpRGetK3e3BvDLWArlRxFAEnqpUI8WV
8H4Ux4IwFrFUyEh5SYNOslZ4ZZPgudZuEo1ywRmAmBDCxsfYm64FlbskzAAU+DwSReqSLCtiMEWC
4PGAws9jDGnk0Lb2YOqSOLvMUw+dwt8dsmbvOpatZ7FLSfSb5bUnO9raXF0oKsS7RDCzP+qd1w+U
yz53TsahXV9OM8iMs7Z8yhMWw0S6hejn+WFqp7yQog5bJkgAg8van0KEhw/fN5bLVbLh2OgMQgnX
XRPJ54wjRLwetSpxJBSs3j5BQM66iYvxM62C4hvigsnt+AQnsRlurxliuxxRtNGlsT1WIh84k6t5
SAECGtufHSlYvttqR0U7f3TAe5B77XNi9w2fFzcRBt4oW2RDpWH5C3DjOdnQEm+SROUtUx6VVfhw
3nvVdK8r5oR8OR078onnK+u8C3KR5J1cG9xscPXFZH1thHu+qpe/lNJxoOYQq3Gax8v3Md2382Ab
8gQYIknuOHdTVdLlIIcp7Ra4BVFc7IyAieZLaWVzT0T7E1hDJNh4J7eEUeB90RktYLU4ZRkc0tAi
R2d2eZq/SggO8OXHj1i0UyhCDdiTNqujoguQmdNHVBvDWmzcDtoBOkdL1SB4686xca7w3yOIMNac
MG6QF1QayY07uo0LxUNmFRmjevrUVpW/W0wEhguVnURnMm6A87aXPiIrL1oh3gVnp9bwkVmMcsIx
Ipg7Pnh7EnNFqHi54IVQJ36JdE+sbq8ge43v5udu/zAzZuniArwrHZ0eQLrPkiwx0e3luOOvvUVb
IJl373HYcwgYiyQ4lQlFsw9m4dbQujP6ZLbv3DcSCv0sfXlH79xeRa6S7IDZUAVHK4E3rFSS3erM
XMkrLekWPcHFYuy3b7r4qfqs22mMxW2A3Z7zGQK9ED2Kkqg5oU/H5q7abSDBKgS1YQGl5gxpHvxR
Vspnv8Xqxe4qBv25gVX8cV63zT4FYQkvl3bXO6tbeVdgMbb0dU12+wsoOyBEEW7E/PXZM+w6spAT
pDwcaiGdPPZ6rdTfuacM3g3eQk11JiI1n92j9px9v9KaAjD6m4d0VcWfWZwZf2eVbHEK8hQFbtP8
1Q34MYIX5x7/49rAbmD/gkahmLmcBB9NbzEzvYXw84r21NR0UHzDN/m6tIHs7iy3IQMZU0jh8nwj
4fH6CNqTyIikXTTYB523RP/rr8+1b1+IN73o3zsY/m50eYGNbC5JmxdBh7U5Rcx4U99xEp42HEv+
bKSz3Ijsxmhhzm7c/XM6WIkDi58EyxkjFcY2uVSN1IYl2kYVb1zzZarE22rC9jwmkkVgw285/iOj
R4WpOuW3cQDTWBv47kxi99/AC1URp/wUOSNnrpaMOcnpj2yUrrNaC8zXba+0SoiMlV5TeVp9Nw7D
m+v4Ilzxt0Qj66j6cGB4QF21iYaf+m8E0wE0lb+7d8U1WdT/5Ob4GyZhpdohKrKHsQlxLo8JJINU
lI8ixAiOVsNoOlyymiS1en2n6YkLaTqjkAG0I5FZpezWDTX/gZ1VjDV6dUUGXnCQ1ev+nUNXQBAH
bguJZwfgZUW97RPyji8T1KnNg0RBuTaL/B05r5n3kShSGTQNGEhZViuLCDoNaxAU2V8U9eDfHgcE
Irrf7Mw7FU4gM4aN2veAEpwAZMqpuYqzE3r8Kl9GaLvCzfxNaZ22Ecteq2nKKv8dxMN7gAP2Rl5P
1LKBcW+5DgaU29Ta872v6UlwOFVmR7Rv1b2cUQQ8RI9ZjzobRX5iZ8m9NLuERVP4HMxyK0lXUqM2
Lpx5iOjW/PakmTPRoENM0lteMe7Zn9ZcpeC5/MusqxeF4f+1pYAdr2Ws09Fm+p1HjNaVWIjlzwJo
B9IsxBeGlj8eRQ/bBi9ilv0fufkwV0XT6eKVLcvOYgvjyGVmXdWIoNcFW9vJ/HCKjH/ouJss/Qg5
5lAMKHfgzmExZaFEyroY5ZMxrxNVZNdQQAdyOms/2sKf15hPOpiFgESF30NOjP92QE/Fwz4UvlIW
BDJcdlJqr6hQh5PntbO0ecezEMIQj5V2PqJUu7clnFpBdV4RxI5GhaDDv4i2EAiCAcEHuguLfHdI
jOnTW6pd5r6qEWJB/dVKJh66hWSRXIKrzYRtCV9lP1+9eLha9F4g++il6/AcQneLOMHnHYCVZhGE
MrdlDjHuSweFQFT5Nqxhvb9G3hfdiodQE8Otlaab8QvOZevSsqpABdIIRDxbWBnxHMZP0bpaoIPD
mUq3N7JoOBfp/BgjtkBm2lepUx3BJhcFOKEkOoT5gwezxRCAMwwr8t3/xp99CCI+0nJFWlSuU1Wq
31oTjiZW3zj5OsVXwQepK34v/3lEiuCNBtpasovXqsLffxG+h4QaOxZ3P5FinKzw4Cg1vusxK50y
5xNj6o0Z5gDpUsI9nFTk/VTxRkuE/JWA9EmFPvYOgluQze1exWah8NPIj6e+K9OluOWTmQ/XmPfu
hV87WVL3rBHdbuHIkcDJz9lCskg1MrChz7vnQeIrKAz/RIl2kXkwQX/3mti+A/svw/8+PB8h54TL
kzabuIuRng92S1zkmilc7rOQFtuhdM5Ts7IL8ulU8wgwWjYY+sv/pboT2274AvCoGZEyNFomQWDH
tegtrHleKt6EjHAemxT7VoC0k0BtBUUZsXG+986+Rm+8scwxV0lyulpmSwvc5tPy4ZpxIVruQRTw
dt3v/1I77lj8EOSz+bWUw3UWaolIiNIWtXDlQdmbETIneZayYh9UijbxzWSmtqXvpjx8CnojdHj9
TYng7lL4HkffTzgYV87l+I3GbSMTv69e1pRTu45I+tnXqmDP6g/Ai3ROIJgsZM/SlAm3fzqZNX2M
gWEdk576GOp51vPuSal9/kX9vPSTg99bgiXh6nWGgaGrqarOyrIwS9Mpc0zrPsnVijwdBTZVMJgB
WonoKBBv1MGCQgY9qSRgoWth+XZK2lR6DVm2qk6GolTXy7WGaoq88NCVZd92pN99EviIQd6y449A
iGXCRuF7ruLWZZWHJjIgFKPjt3Uf2piKf2Z0UNZqd3t6/XfjocayziSYhZ60/YpOtC87EiEOJqY+
AXQaxVZM9V3lwEpNkSCNDSh5p4CmWXHDURSR9hm7VPItjRaFpyhdkgzspOvWSGGe+nYmAxtid+Lv
9hhcrPXFxezKZDpNxnHf/Lim6ijTSJ+R4vpaRf2OZ7rLes98MIsQOd46QbElHiZ9kgjbJ2lBUW5O
zI4c8GTGPcPHrcdTndbHpi7lL+Mo9hWn1e0j/AWhNJk5MgcDJEeT5wjECeSwklplO1U44uNtamYB
IZ+gKRN/dT4AIrDoLqvvi35KBQMWMQYtaqHBlEmYQGQMH3xozJqNH/KbmyOu9TbmOZos6INWM2we
4ppw+4WvmPiZHS/WReCJtQszlKERJBJJ3IqK1cvp0Byje/w8AmSxrnP7BThFck1nr5/03ZYzFAdX
Gza15D0AG8okrpkVF827hqG1qk00BMopQf4tB6T0lgBNCA7QF3MqnC/iWJaB/t6VkxKgXMe0oWki
LgtaNMZ5oD9c25oBdw3m3O30uPbwzIzPfYuB1NhgNLL0mSSA+o3pSjw835b5jDAMw14bjegO9bYV
kvLuAfeJ+Hqmj2iubSwlDgR2hIRIZqDn65u54lthEzL+RN/VlMEnW1dv6rAXrvq4tqFtMlqWs+F/
xUb1OaH9MFYfKmYOIQ0QwfHl9IJtj1Uq+wY4rfjWhJNE/9Y4+3VDRBe+gRgMfXkZhs+jPsQNKwUy
oaXIHldsNmJc+5B8Xx/+g8YdChecfSjDl3qTPYeDrCZj77Pmvn0sXmmQ+taUg17G8Q9VAq2x1O+1
Z+jJszE4XE0yiN8K4+XHs8tE3fc8Dm4EOnqupuzZM7/nWECj9dnLPDoKTvqrm7kHdhiiYMAr+0Nm
bgl3sVzFMokrYYrcqWKAaOkt3gQIXa6/G8Usp9cMdN/g/GNNbuMf0t2G62Lxn527Qv9pmHezt+B7
suUyur6FEQ2ky5QcImxYeZB06YE6V/yWmnjQ2TXIm9zTJao0jdlZI/gGilWLUxeJYWxcjvAZFWxg
AvPyfVQs9tJCj4U0O+gj7BtSUhD3hae7Rb/legJ8hRA1JH21z1oTXi9h0MaCkIZx83P+2IW+1x7W
SYJvyZIO5CwyVZO7/hUk5293DeNw/3w+raT5hJcjikfK2Be3LlIf5QONTsPX3MRnfFqmxiqCQnJi
qPxuMA2pn1FhEnaFF4+3bWF/xwx7r7Ux+0rP5OvNcEpv9R4Mg7oiN5ax/NtmxHICmX829YLWxvfp
/y2qjAM+4WASiZQ1oqi8RFFwKuTVGkWdBBeDvaL1kMKCOp08aQ45cc29SeOFnsvEFIUEfEkxC8+/
sit0+ukRgTxp0npQDPwr3X5OG4TjJRUzTAMGPVqMRvXnbqL0+7PieCexmcO7mCJ1HSlFW1nU2shU
PqhJL/jhvMaVQAmQt5poT+irSds+0/320pBuzt/+zEFzoqOFvGX/6AQ5i3ZeEztsYuoGwFOHbZHd
alHEDoC2/UXcyq6dUxMtbXr6ImA1ACHcWZbPj70GJKcInb+Uf1do1Phb1miDwyTJYV/zNDALZFaP
o6JuhdLQWFCMzA3I+G3QbWaGHsJaARO3YNd4jC+28mzgbwxxQx3SahXJ0TifjTpjMLIzFvjrH5cx
f/dZS/deYxbWyo4yNY0sLsOCZl8HURrf1rATjV7++AjbkOZEmVbFlF9oxUCjBdeCEfxjyLXywDOg
WOKC4rO2I7gNMG9XNJGs7elS2YqvCsLLqQeuYb7/G6X/jLoANuycNLnfRBJYBdZ145w7ioLcNXgy
ma7XuAcWwctPJg0STrutFyzy2LuqT73HprCHg1Zx8QwdZS0xdd+YRI7McDaO9p7wMC0ubqsAN3j+
YJZv0IBpOuqOZb7LmeZArbIWNW581fg9sf+iqwLGmZFU4AaFdw+lz6sSiqB8sw4S2JmHI+FWRd2B
vAeLNciwEvt4Z6ScCtXV1EvTV2J425DhkX8ZOy3+coR7ri5vLmz0zVElqQfAzr6Fq9B6U4xbERzw
nCovvhtw0L0JhRkWdIBxMbNrYTi/iYmQKfBwLgvJB+kx5hLEPOmo03YpBC1ETKPda+dTt9As2xLw
KOaSIyd9O237dwhq5WMzrHBN1xwtN46H5zNEbUDJxqQbTspixP7kj+cFFNHiPAc3ng49SzbMJy9m
BsTUoXHhPnxEXGs6H6mGvuRwfyGwdWbnvKoJlCEbAhwWTzrBOeLirIQbJjOstA+iPIVgDGGhXKPZ
JOSSYAPBTaaFAhue3dvqfzJVPYbX44FtWTCKsbfkl9CreOkyZxuj+Op2LyOJWtnP39OYgzLvoOYw
ZI7Z7gcTUAJMJ0aO4O9tlS8jt8WB+fyRYWF9B+KUxmiTrunrTSA9Gg5aehIc0ZVhugDQK/KxWBbr
GRvHG27PO/UR+CSjznr27IBZ0dx64N5SPUjddzPyGmH77HPhsQIzrY8XR4z5/hnFQEp6WOQwfN+E
IgIso1FUB8qy3zkAKEcv17I2AYaXkfrhTgQgm2L/BXY8z2o50XYIJXnU7hpFrjtgPjEdZ+3oiF2C
D9JlhuabNDK8XlbQ10HlMJPX4BhwlXvuSwYYxlGURMOIJKcqNxAi1REdNekYYEUzF9wTll2dFlD7
zk+nkDTRrtDIvFY3TFK/5c0QbQgEqPilRggWZdsG+Lv7ftTbDqyYTWkBKBuCdG9W/T1D1Oxx/g7h
JmWIqGI4CH34d9kTJ3fNAe+sJFxWTNgP8uY9c+29pKhh2NwlmkAMHHS9uBHWxXxpke6KB7qhY8ZF
pxHHvV0k23fHfm/GMtGMK5sWzSCYBQwDbHqQF3TpNNJnqjm/bwAcmzCIrtJgoY5fKPW8TV/ctbcQ
lcK9TjOr/dIat+9/oH+1wL3GjhlCG+dT+dUR4I57U5iGAy0ICZ25WDdk7e/ktpSx5GMcw7oTIDLo
zSPHyyDd50EDYBzvONlH9JfewcPg5mo38XN7sRWws78fA+0JX1FSBQNn0C4gramg3EXoOoTn3/Zi
T6s2LqvBz5FGKskDTGVzH+8Ommm6Ab7TnTEM+STOkKJjehiJxmJoLx6fqQ6sREWga7qNmunLam2z
l/IbSP0zkE9AIlbs4VXecSdQVySMife7L/ezKV2HohGIDWoPlzEpsLrCk61a0irqbxVvxwhfOFFZ
WWCdSsQAYDGKTWQs9CGCPWsBdaQbL58p9TppqL/q31r+iUbvHMKaqhNOGM4eLdJDFGy3MBDTxxs2
/8MVAJvzRrhx+qHGtXxHVsewt07DTxMf0RMp6FSdYG8POK6O1r1ibwWA4xdd33zVsBunKCEeue5N
19uGEjhImCrzdIDCDtXRcJ8M2+f4KMDGh+t2MFkz9HKNmKqSioLF7t8Xm4UFgbpyaUfh1g/Uva4Z
i+XSFXAWby/G1CzeED9L7TYC5q4/eFDRhgQoG7ATSvbdkIuSP4I3GLIBdF9egXtQE6RtIZ3VShNP
6s9IFJS/xtuUK9WLpRYqkGUtlQGC5u99WxX2lRYGtGYoCiz4tFq3m+0VVyjeLOa//Vl+lczYtmv5
/Cclhi56X9bjVzJ9kGC3UtGSPu50RJpxm0fvJOt0x0MfE6a9Ml0EDJTzQb4hAFbWyuJP9WDfOfBi
IuQfD1aejhLEbq3U6NUblpwJUkLhRR42vqvPWWmQaKVYq0wagU51thm67WSOu9I0LuBFqqmOiNYk
XjclrAN544eGBmaGbz9gqD+uaARgVOc6iCtBPsZjVTHSHLpRNL8IN6ZvesuePpwCop9ppbHOeozh
X6gzvf9qwdPtH9GaYXciheatSX8qKxD05Fv5erRz81XZKnk5tTw1TqCN2TXpS3+iGfA30lexH/bM
7AGSExFaPXjX0Z9sR22uNqsA4M08CvMpB4VYha5W4w0cgM6aOSPcZxZ25jw2MWwUrB3Dz8p6fvuq
srwVXMT8RsO5XFnrq5Y7en5Q2Qwp3n6cfn/PxYCUiLJLc9gfcRpjOW2SEan87PzS64Nj0NXa87r5
P5u3J9Y01VpuSPIuI7EFV7jvznoIv0U+oipN7zZfs20/FSYrKvq+cxDKnUtZS2wRmt9/wLqXkZU5
g8Mvm05coDVf8E2r11e0Lr6c9Qjgq5WuCTjoqBh6FMF8dA0VWFqBzUvLcShyaH3twD3XLXpQ7Loq
yqHrIHKTgrzgWnQrpJjujJUbiFyX7mWVFHtIrX0FkCyarZufqUH5XnIPLd7JtodqurXCI5cxhh05
uiGgCqVhdgCxIMGiNIORJl9tWi26VjCLb+YY0PR8XGmrFMGyrCrM+oPYTkY9SyiJplXGs+gHgHrc
8gOzh9ZAWzAlSPYjIYlESigm87ORL25S8l3C25dzWLYxBPdY0RbJ07YWqT/HrqhkJmXyo6D/CZ/R
bWuXXGNXWoVw8gDs4ElvyBtt6DtJCdbPhFy4FUguziqVoCDTzFWvU2oDQBPSICiB6GNirT5m9tmk
KyqXKHJ7xubRqwmEUq3JmbNh4iJTqk/SmyyqqLSJksiukMBaJ9SxjDG7MPACjKhItI9iQQW7Zkyg
Jhl8H3gN84dpKstSnsG0PJm4L5wgH6MIsyJy42TkrHyW1T3Ap6cuvpgIhgsDL+DaWdvFohWzhMgP
H4wzM6wwn5V/6GuFo1Pmvy2Jw/8LcAdsV60UHsWrBzJ9T1YzwQtiMk3JDHR5YvUMJOADy1I/ZaSA
GHRY8LJ4XngVdXw7/rk+RPDD2MiViLUwqtOFKfBBcSlVAHXHjSsRARo42kgIY/H04SjBF1GmGEhZ
QrRk4pGwKRXz5KTxrMNy/gP32suOlDP6fboTP68BGtUpOnTVN28poxW1qp6mCkI0puUJZzbYF1Zd
y2rpqcmyVwzq75VVrW/AtqKUqUydey4ybqPLPwE150npK7VLSWbxfAf+vF07anC2Ly1zISc2GHSz
wBLwmsKiU4zo7NxnhZU+UGOz4CE+RsXZE4cda6+lYs/AsdNUKCHKuUhs+pxC9tqpHm6n8KwmzajZ
zdyjRMGdM7fd8GEdthmvxzZvsc9+IuFTbvhKjutjaXSbq+Tfx0hBzmrlreAFOzXwPNy5JDcoimn9
V+B9p6chJmGqG3DlXwL62sPVHMPwWMSZGwYLAlQESYsuDGVLQOyNwCoc60XZ6uwlxj+Rkkg6ic55
3xOzwwcepK9DUrf7Q9tHyG34+xXfA83RRTLQ+ZAAKtuCxgv1EMQzPBnYk1HkfTvTvm8vXDeI85My
t3hizB88yypEKmjLpVudNhZraTYthNpGV7BYxB0mRrCcDPV5asD/CMSL/UMzPCyOQBybPvAPrAOM
xgyhR0wgMZ8rPmFmi04UBBgKHfTU77wMOx8m5oHXWON3GtX0zCbaWCZEVAib30Ciw9zSdECPNRTJ
KODbDsNK8oiwbIIIba4bqbFaWFm+LBprb1PFVGugzghI2Eaz2wtKTgLkOtsBdwTxxxTdXPp4GQpi
zLrp6EI9+znHtDsBnEtmg0BvlVQyhLT2ZNRjL16UFmR35MPI6FPGmMnNV5OU+bJK3iXdhtXwj4lI
XFzjzk5Sq9nWPgm2OTU17wjbjAxhVq3bR9tb5d0EGas4ESwWej1GxvL9QWYwOLvak9/VZgSBunov
RTeuZtGt1JBR4SPcaY5kinkcCkzbeFl08sf7y/nc8T6ZoF7ucnYqJ5vAkWt3Il/t/i0hP8Ef8+JA
DH1EYdk74Lbg0+CH7hc8TZ8adfFmM959vu2tmU1jwhv9zmeNAQ7Dgg8t3EdUF7l5EEAiJIdlUcvm
ltJ3seqjCiWoEv5vFEk1sOc5+HfVV2nBPiUdIxzvcW6VT1zCuurHNscXaIrHHw6xWiyVkRFQRg1P
bgVK9qHkNw5kbCfL47LRHHYqaDRWT+lSQkALu+uJTGTeuRU3Ub9SC881v9O/pCOskwao0MG6EB0e
lrRvPDIQ/tBsb9NUSH0rchoak/Q8Sm4W20+FCUSBIpTy/3F6sv/C31VXOL3lJ7RSyQe1zediqy46
cG7Ud2XG5pkEdafArGevoK2QQJuKoQHP+ezpDE2OzQtn+yT5cKenfXaYwX9zFYv/Mz//VshjmJl9
9xIvQqivvZ4GiE+TpyFdMPxqXyMrkmMme0tT6iRsEtZZG3NLbfBobxKOBGEAaNkMfTGAX/ukgN1F
ebY1H/9TwV3UAzNrG8+7s2nucYKsI1aC2rywagt8wfff9wWVl2vOIiNLkHotKPocclHEs0FfhPw3
JLt7WHB75sC5eCPDNos+LRCiEIZdatdWEA5fPZ7v+pNugkN/+m5PAI1VjeEUT8k7n6wpTkESLR++
20hIaIIC4DMBjALWNqxWspk6RV2mQMESYxhovrEVemZwyWcYcibW2yYERSO8v3pVDxCx2xn9y8hL
Mc2e0plfzL+NfdYoZtSmokFRichpfvrdYBHNMfz0Xr0hWHFgAFu+188TuIt1dRUxpUM43lf9VE5s
KLv/+P/pk7mjpbM5g9wFW0nvZKFHJDAQVELji5jGgiSxp6YtV/9oeT8KNcZWa7XIOEv/NZnMNbHI
IIvR2Sz8+yXfQtCO50JB+x18w2fi9FYYuee33f3A6sPQkbSSKlW9D111Bg0yzlCNqZBz4FZL1eJR
1qnedO9OpAtic9Bu9BQajhd8rlKttuCJDKSJ4j6h2nIZGtmHFzlze3Y8OW/2g5JBhPTlKvjPnop6
u/KcnwDO8fOfqXYYdwzZ3hoh1RtoHqUVbJ5PLnzeCB5P42VrFp00ZDlMcHH3iHBmR9ihvcwm5siX
6vinlY+FfLCCa/r+ucD4Genm8fSlZN7O/u/9/YUfW0tYe3/9QDk2v8BDk6E7J3AzYzW9uzBqWGzG
PThnOZx5RuysY1TrXbLYmjVUpKwDQSyjvueZbFu0KPKJQ5ORukxd1rAF5fY7g0yvXR2EhZCDGLfH
yWDHrHGFbii6aQGwgHePdhkHoIKX701gN4apqDGF9/KyWHXgYNzQUH19ywCuczQE+Zp0FRfnf1SV
ghQqN4tvIyB0CCoZFxDKEr8YpTwyUAH497/E3IXhr583fJvPG81z3CTze3UTx5QWffvIwr84X9D9
tdIgToR36KrFn1cTnSkN8OBTxqNDn5hVUPjZ8zTQaPjJZVhP7uOeKL/skoox1tpkDYONAlfs7S3r
tqzE7ortGjKBpZ8KhMNrOtWui36chRTH0KAN8LTJGtaw3PlaUHtFjEr0vBitCvuB2ggjxSQGMKLo
/SGyI7YlxCQzbUvWCwCiiVRKzQPTulDCCgekP4CkbAm433+qjNjAWDSi278iiaRSwWR+IQXIs2Yj
viwCgsJWPb+r2yRVt0k61vLuvtWznKh9SIwkMEWv60J3x6DvqXEeIBqlJzS2yhlRP9Q1Y+81AsHv
OglR6QYOzu3g/cF/FqwAw1Eddu0m3Ki53Riyl2y0lU9BpWK8E5PODWsxkGlUkCihx4+URv8gbfkd
PJlwW+oppE6fkxRUCTc9a6rUvIy2C6NdiuKu2AexNhkfUL0FUYn59aENQArabgeo5AzQFQZkJFJ8
HIQ9nEaXSJ0kvjDyblEKl4cfJcIGLpjKjxchFa/HKcA94/jdSP1PLtJqeeC1QpkaC8Gexymv/BRo
XajFNA0++bNWJohpQVcWqk5RHOzXOorrLzunr1l0zGjmSt9JzxKYrRBTifXyGm72+kBvGCFMk1p2
bI/ZVgfG/xZ8j4pYCgjMKR4VuikNAdtkc+unXfMBObf7aNX+Wz1FQMPn8dqtoh69fEXAQu5TCpsm
/UDeGh3i2pYurMQBMyv5mAgjmDPhNXysluOjRWb6wpufP1Bje2Alby6sotr1D3Sl7Ml+r1Doo/tx
8OObddtAE7qrdMMU6Z4jWCGD9YuVGBtbCZFq1gVOLHMG4L/FPXz0CT5wUxP0U0CSdCaaL3ssosAR
SmBjfaR7eNLyidTx1Eag/oCKTPMSmcdOl6QkGu91kcNrOxqZJowBW4JVl7+MEu+3qeoOo+nF6/pB
l4vZi8Q6WLOINHwo90u3s9IO/wn+RG9bi9ey/Qrk+o5Rys+p60hvLQu0j5jA7pSCB2cfIfTlumpe
xg1tclbzyszorlnGkIsbv4+ZaT+s6OvrdBfC9BwD954wWYEN6o8u/3xdRakqM67tYasQ/jK0RSCI
CnviRr1O1qAAE2LKimrcaD0LkBoBU++gaXva70rqkiLZWyNVpKyxxB7EkHl8u32HsPPeqydJnTy2
oCUiJ0fDV+SyEQUMikH2Bo0Oiiig8MlOS990FY62hj5vsu7ytPc5xAqRSwtCuyJ9XbWMxO1xqRfw
uvCzYmJDb4DdbHQnBiS+ti00W428LRqAI8XLUNYlwBrIan4L5HqwyXsKIphZFmg7aRGzNxkYRGzE
d27k/x0+dLUWuQio7WVWzcpz6UYbdS5PYmHRjkYC0hA8TGkUDGvYX0Vt4PA3stxXXUh6GLMW/Rf9
oO4KJXhSf4oPBTisLEaeNRME+BGWzRH4TG+GkP//zPig9pp5XSbUit/EWCZJFD2PG0xoZ/m7mfvx
ed5crFr/npLkgK8r1YH0vEv1lYG2ZXho2VGy/2f5Y7en+mInXelJceOQZdwggCkIK/uxNYpiw65R
gxa0Ev3z17ePpE4E2pIuP+TLAFWvNjech7s2kfal6bd9JRlv8ug/DaDSEbnhQUPsarFb48hna7pV
wXaGPeeOANgz8B1lSrLlgd2EHSwXAK+C/e5pKa339yoM+Wjxoczlm2eeNjL27Ht98uC3fKgeIlCz
GIpAgO3D34DEK531mXCSlS0WKyEKc6NvBHGB4t1DCOb+9Cb5kFOTZDcnFKDrJqbI3k3c8uomdYfA
wc35MDM92ZZfKJ+/1AMtfJoZsRUMu7zibJPij32jsMvlURtj6u7Imhbrz0wg9QcQvzw2zciJhIcR
WxnpslOQb/GNXqImQgmncKisxj0IA3kdSsuIZwO6i4wGyQEhhLBDsCtagQ/zR8ScX2gs3egf8Jm0
iPPaKL/lqmiVlPhxDvnRO5tm82g1UuM0KXl88/Cb38kHFxk8F0320vIVDcf2hcMPNYJLSNErQG2Y
s1/QrPVp+LCC201DaPYkOTufoDpFm2QV2LCIlIN27AN6kc3I6zM/gSZYnNs7fwJpzRRPVzSPjIm1
Q2EuLMQCy3ZGTonRmPJFR1o8XY52Ir334y+Z98OToCaTdLqY/Tc5sLOmT20uCoOpI4wkKIq7jL0Q
HWdfOdJl5Yqrb7HV00Y5tdggkHMysPbmrjzIYn1iesBnLnwytR222Y9/HMYZyK+lObdjNkoaCzys
2fpHntBzSxEYkDnWSSaHtIPg7hxXDfeHwGm7dhMDXNXLJRzckOAspY23MZitsKTXzWW0X2RNXzSY
3Qrtnr442+kd0iJWtDjGC8EoGSMaQguo4+0gD0VpCNmn2qC9M6VnvEOVea3PUea3+WO7+RyZdGww
Sz2met8D+m8/q2FmY/SyvgjttzsTRdAIqzua3zIgwz2Eu4KkggCC8a3NpxQ4hvqbGfYFZJO+LNUq
NtqMGhx8xCqy6YFnPBt94wWDCzIUqD1HiVuzEWnghAZX53NnILvycBBlReZFwr1ChjYCB+cawETR
Ejp/JSxcMypoLxaDg2HsWqXfVi8z9QD2dCpTCxqhj4UtcKgFcraGEBI6uJ/ss8ym2ygpEctTKJs5
ed8ZRPm1zh8QmGXdxlgF6JTQuO50K6KdkHhjfOpHO+3YAyp1g8j8YK/9WI0x1+Hn3p0wpJUzURP2
vZmwW34LSmJcvukMABeWsrQJNJu98pT119MsfPpnFHBt8LVFuaLlO2WSs4Ai/FtEIUIuqqTiK7up
cLVNGLtYbiQ7EAhS08MypEx6vLRr3xt5dDMUKKZc3wv42+w+rrtqmJQOxhzuge9XDODeBTZ/c7Jg
Juvx1EFQFzvY0PinrWEF5K8wFZaPkuc2KFHHlEbwpe8kwZKayq49RoprnhNGoxtwuBIMs946YkyQ
U+/S4KkU2b2LY7yaUSqu8M0z+nMJRRS0aVXN4fB8cqc5+K2Nb+Um0xDvOvS26m36SZvgpDRZPMqk
dy17uV4xifG2yXVLpAqGKt18mH72UfnO9SuST1yP7aDbsY4YOR/nvYfWKqpHVwmT909dEMaV4HiZ
2kH3bl6QKSCTph57VzPHdcaAZmHSVLTPW+Xajl5whCHS5L7+eRRJImJveVEQt0L82tF0tCoithOv
Zm7TmWDajR1OOE7NzeyGcvjVpFImskzeegKewYnj9A0iWfuXxJnWsZcu+Voun+DBhECRnO1dS8sx
ZeVmu7pm7g1JXdw+6JM0yH7z934c9n/nlXUI4+Iwj6Z2lzCBniU60uGR0k7cg0G3TKPGuQnN6ymb
6dbsCop7O4h4MqyxlZGL/ykS4YrZD4qd8QlCt5CurTlH6TgsyAvO4yrBGHtx/z4/bn3fF6cJUM5y
XX1rYszRYH2XAdWoq9X8zQWZ9VN/yTkW+eyLYzp/VirJg3x4Z2zJcGNlCK9zoSNX+7UNKCXAgcuI
eX5TSK1Jluateg57zv57YgaVP0ZzPO07bVVb2MwCYhnz3jwaQzllB5a1WLEpU4IRouRI9+OPckcG
e7WedaLAChSFMmEOy4lbom9YRmIRCiBtxAv7i1uMNCVi9Z96tCfOwaVJiZd2tOL7isYJI5LFVWZV
XDoYHjka4XPIOKmBIYN+Y6aG4eKXHS74N/Mo3Sdr/jKN4cDM5FZmTQeqAhieHHEGr+mgyEXGBPdI
e+XY5SbFpNU14T8N6tyK18vq2mIoiQjv1cUWjIf/yQfvzW0CseVzYVJovmXuJniU1qn3epPDsZZv
ZcS66PG8oKBR1L3nzrBtbsOY4S5O14fHtwb/sBzj8b9RNoB++bLMSsoFvBVy4t5Xqc9HQTjWV7fr
mSU0HCbm4YXi7Sa6fr+l/fang7uOQbReODmwKKbmAOnsLRyFsS2aptoEGp0fLclKNRl7WBi/sLIr
reA8v+69AX/fxAdU+gWeKPVS2Ztf0p+Owy3oei+QbfhFac7yCGVDFq46+L9ulHY4G8s/ja68Xe4y
L16abTsaMoQU4PEBl6vw6jvGqlXRnMnc0dl7xLNk0MUXcRxNKTbEf7OYfwuXcCeYnvnG6Uy0GrhN
yNsbPrpNtrY4cA18BwIlsFOXc2KM4G1Wu5hRimY6mNHhyvFLTL1pUJwD+A6TzXtKUQC8v+753nlw
EcFKBF6hJwve+MQZcKnxJN2t5JItpV63tG5knz+qsmeXw9d/q31RivTkfhm3vWXZdPvuPlCp5q3M
JOKC25dx3hFg+4IdEHXsguxE7TrGpjd2eCBDjk7yphdcGiZDVe1xwvLpBA8A3fXBZd+SnhQ97OWE
OL5dwuTBGNr5oquMIdrvfIFb9tZ2IXNKHeXrehxnM5S5WYbwVHv7A0yTRjcZ7a+6F/uUb31wODWS
AGzOawpRnFEGEVCH/k4EjF8yZgSfgDlNzKxq/dvRl0QByraKy2PuSbEOPcp8AK4LQT49DDw1pJCR
t6759UF3bCOMlx1i7kfBLDhSOxaLf2Ofd9BwllgGcK8sz3ZzUGPs69Gx7VCQvhQIKZnHx9y6PUa4
2+YgOWnQekywUHVyjbYdM1Ph7TDXOUhF/6xQjdIPKqWqUjwWXbkv59gFdl71mX9r56xTzPftH2pr
tojx0UqHlGgrta5vlrf+QOFTDvNQq2u0KeSAu2Mc/X/nS3EbLSvvRbDvCXBg2SQj6gkY49SsoQrZ
MBrvCES/Fiu9cZ2e6k2bnG9J3vmiCF+WBDOaD9JKiiSMRQyJW7rOYjr9WNWYUAbYKOuSiiAnYUHl
Gv0p4GoYoyCaBOlhydW0uWaI1/7yYjcxfL0/IiQ+//Mr2CwtYpJx+TiSIUxPaw4zNf7s52PTIRAM
dtaCrxxMjYGYUfmElLivLOgO/ynxcSDseAGcxEH9zN6X3ajGGKDjPLSxgnxsmYEsaev3rCiooIht
te+w1/NIow/S5PS2Qd9U/TGaBZpd+SQb6OxyCdoJVVV527CqNLXTFqRhH8oMM+OkfgvDiJroZWMf
s5/ThcgxXRZ9hm1cPcSu8zba2KXyca3OivhUeaZHNrsQoCgaj6yUhQtUl+G+ftDZ9FFSQxl7rNx5
0pTgP4nTd7adYGPtewqgxRkM69wW+JkQaVtpUYt6wadztY2JdVZdSw41uGkAyWAa+SJjEJ7gmIRx
zU65zYCjuEIvza6WZzYqDLEGwSiuSi7tpC1XdMbhKs3nAD9TCvO47ulrP8D9CKH+m59EemA3UXSq
qDQZKGFmLXi63ZRYwa8rnQQZIcPlk29hWppFxGk6uZFi44VxuPxcVEl9kcerdV7g0ZjnyjR7jPjG
RCieRGw4A114lMNvU6uN3lfdkAK2fKRv7Je5j9TsPcmGOUAW5nsOFIkCoDyoBHBuFJ7s6cRtdNpV
LtNwvpDsqOGEEDHPnJSHmUX9ML1UEhoLgfE1/lZ3wg3cS0XB3LefFaV1SgEXLZeq8WpVQHEnYDmt
N7FlYSIuGPw1RkVytyA0M6Dyt92ApOWMU+6Qcvk7jQfE25cX/cAT8LyieOzsYXVnUFwsYtnnSszo
SqB3FbK6d+MzeWCUh2MhkKMZLQ3VmbNDeXDBoBbqepleni3v7dX1TruRS3fXsZ+z0jrGAmiOqkXy
mwiyECBDt2ff0JCudMbT7rAwCj/ktsk9DVvRDrJGNIAa3f7euNP6unxnY8Z1HS3obHLcF1ENHJe4
WuGkNwBZbMDMk2qtfEkIyqfUbMRiChhhK7Agwx0yJ5bx592cWBJlG44taKYE5OsP5ZiodHm3YqHa
gA/byGEIkoSINtNRjzxn2L+BhvIa5n/w/gK42Hg3CL6N7HkYIZOZMbsMQSoOEoylblud9VZPgbno
zsfyb2iSdcNg27nt7ReuWmCy7vf7MAZac9S39ew5Ti0pC0BQsbWV+TyizWg97+CFWY7N/b5jkSoL
AW1+vYz1toMwxVd/+fSeLVhtYkki6FdD4OI9oS9t4j8tFSNQCq40S8zW2mUQEuVH1XIBBzIDlH5A
fbeZewzks+dfNyR9D4i13MlKo9OrkYqxvWZrpedLGOIheUWdLnRcc+ZmUMhcq3zW8xyvw5ilg2hf
VVS9YLNT/PziGXIKmpiv0NdQobKpPx48jDq8QDpvp3pc41gakSZ52y76SrXpLM0Ic4Cw/qfmbv5m
xOUWTHDqREqg97shcAUiibxzoIbzHk/ewXj4SEY+S7ZdWUUt35Bj7KWG/LDMqFMGN23GnCH/6ao0
r0b7i0gYNlhC7YYhwDEhRabi+rm/m3sZTXK+b1NfTQfU4nfuOI59L0o4epcxtyd7J4j5Nt9iK6uf
YzYU8DK70W5YtXsSfta90wyJEM3PFbCuaeuxj1tivkM3h5ByssTmrjy1ROw1BVW2YMnGS+yfxmVP
hsbTN2kisTHt/6lthmKMfUkL/k61Ncs/qlh6EF3e80gRhuB1hq2Be6WlDEg/lWYaJkMAEqJkL6eg
1+TH76f67ceiOF0fJLnRgwhhKMlpdeaFoSbBs4baqRGMTG1ujcWij1b65c6qFt/1Q+iwGKnnWjs8
8n0X86qgDjakYYar5wpmN4wUMJprxFV8iXbn/e7IPbveLmR7r07pXCdrSfUKqycY4yizYHdW5GJo
Az/WRKnl3TwlVub4T2cDbtRH+1SrBfZ0IKjXi+W4zCG9yZcsk2Ki7WilT75TgIMxAw7ANQd9QrEd
p3mwf9gnqMjrz1vBx2p6Kh1jTHfXxeAFb29E22AqGU57mL+PPPN0c9daGdX9tHg7pPGSgr1PT+bR
Ft8OYs5Oqxz1ZYxEYuq7ZQkuVeJ+LknWZq1NbNKoQ+4R6PEYUDSVHsJFSBpiKqkjee+zAF0ijZsf
5oJbe371qnZwMMY/7KCAljflcYFJxP/C+RT+yqw4ldmbSkWXSq8FViSlzBcmbNhgq4thLZrXAZdq
5bpcv8fTY29M5PYjy8F+XpAEGkyibhEv/+/qwrriAEfq0mNMNHW6tD3S9Ftjatks62iNhIIIHrbQ
DV8XDXmKX87dHUjiOxtDvXY7h9lPyCRx3QfFz5H2dPFA93cwa/cgLTZN7Xgj3AOWLqeN0Ar9PTAS
sHXrXLE7ymSMW3Cm+1EYDoUwxsSc+tvgOmEwgvjwZFT7bdSapblleB1+lUdLWDOUr980ktvV9OmM
3D3x7U8tFU6PJKODsXf14wa3P5NoFradppeEaNY8P8rxzoAhXkUNq/sltGzFL0sM8DUOj5bGo9Mb
tEz4adENMkUkATy6j7FgHlIXeRrY6+2C4bZYdIY7rgsBa8Wg1ZQYapeQ5J6lTTjxSv9WvkUWphMu
m40z8hUROwi6q9P6+Elst6axPGmhn8n3NSDN0TxWgU2isyoYmvI+tooYIvwhAlZV6Triatiar1p1
35twL+3IIv3tThEUS2rSB41fff3HV8DEYE3Rw3MLFv1GdHh2d/OIRmKpMWikeXKd+iF7B5AMPRmM
rQHpmtmPdWM5QMsd5uY5gFFiRZo04gcVMfKo46nwaFUcB9eU8zBVSFY2opCweANKp0KZOVvQEj8U
663m+neldc5xLiOs2cHqcZzK3imdBzf4n9sKymN4GWbfSrWOotGZeyhiLt3ZOz08xSLflVR4ryLf
/mAu6YFt06bCqRJPMcfvjktw2RKx5niVSuF5cgtJQa6WqwqnNkYdUymGe0JdW+PxHomBI0//I+Lq
gQSrob4BQpaDBfT6wQEqEq1wO0vgPZh7eF+IRGi/KKm3x030w0YVv54LK4TbquJ3ngZo40h9LLJb
Vpbpg9Dr9E3fOCex8TvKXccyAz8W9yYE3WuqgPf/Wr+X5A6jTDixUPolhGYLSslQ7e2mBeDriEtP
cZqmlKgqBAJEYZZ6pTEcLu7vnmLdtZNk4tD+kcpfWk1ZVMxIM+r1rBJ754kNHVySpD83ScDGKP8N
zZVgrHWEDVyd0dpjLF8MGDRk9pqUEp10q6XZicAdqEBATiuwxdUlHJutqcgiw57svWs7Vtn4lGfj
F0pjQNyOMh785aGFuZjTRKH7ubWIi4ZbEyz+GJxuCMAznFz9wljQ6MYsW4i0WWYQVkh3NU9ZHfmO
J2aSsrjYtIQPk7Psbj1KHRcGQntv8jtwQULUCHDDeO9y7qYEiz26m9SMuZdwmAGmQn04N6kAZaQE
TSSDGOfYHBplQjxOdpODvPlt8W00sLt4q+9YXuzZPn4L6G3zb/21L1O9tCkbwH23gqTaOXHJWy8c
HlcipmqRzDL0LMgQeve7aErK26z8ZG8P8W9pu7D0aCRBc9dFOA8I04Ur03OcsYO1erzySNN/NBIc
rtoZ1u5w73fQdf4TMSxm5CnPD+mpAtmFliDqk38jU9qYnVE+4hlnR0LG3IXTd3zzAV4jXyAzg3mU
5vhS7oYP2bBXMXLKtXcixbRb91XGd6OZkmCeGcMnTQqxrJBs0oZ0wgw7qjuRj8ObDNpF/XZdvKLU
2bDF2ydbW7Y6Bc2gDo7tYn5S89ZiT917YhRxxPUfvTuqt5pU2uABB+jLbyMlJX9tOntWxTx+hoa7
a9VOlD0wDGq0qQXdiZ5JTwSkkSnGYg4S9wrSTDZiulk3tPU5bBog2pg0U31DJ67T9tyNqdhmVTHr
9H22ZLNJGE6zivSy6aJ1nroqlcjAj4YR3qQCVMgb/mik5b9PjmLvEUcnVEfe/5/teUj3vJfEFSsh
Dj/+YklBaieF7Y3MvVFFnY4cyjxpy+wThE2wYTj+0aRXm8nogBRFh7tD2Ty+iskNOQmoTCmFD3cO
mMrsn98z2YeS0xSlEwzBwnWykg9qdi6JD6BY9tk/27hzVLf7RrFgGmwiPls/hR0Wtt31JiMBssdS
9jNodCmTHKWKT9x5JXCCIXzf+Zmf26loV0NOOEW3vv9aJKtQxJHB7dmUa737p7FRlzBCFnodDaC3
dcSqCkMlIsv0VO/sruIIKQajFmcxZppiKWwaaXUzEMazJb7yN1o/XCKiIjbgIdXuCzw4xo/6y7ko
4pH2M4GeyN/Wjd3FXy0T6MSusRKKwhRI3lPjTylqtH9SZ/vXbQCjCL12NKLgeNt16iC92In+7yIT
Lib2VsVdatc5u464DlAeChBUKHqfzw6lEKdd2ieANZxbvZlbCeJ9k50bF0NcucPusgtffGmOwAi/
myeDMeezqxuhFhjt9/XBEspD/X16Agr9rQjaVNg/ezRimVzXbxlft5mykdPhG9XSMYqFxj6IxGG1
QRnClF61SFj8I9ZYGUiBgkPs164sucuuCABFiKvDtjXjuSmiGUMTCQasksCx6Eu+cfKIxDYcxggh
PjEpAPUyBQgaPNOjqCL64tm4m8JHVQWHxkWjqS9IbwLPCKgFi5ngUoqK0fZifsmELJ7NfZKIV3lH
lfs/4ll/hlzm3ggyAg1sN3FM0Pha3zS8REPOelt+CtQiBFjwWnHIboegZ29fN9NF+R14CfF9WgnC
50HjzguHivTdeFJ/MJjlYdlh6ORuICkhv1gnkeRo+C5SESKBjXoWHt4tJdCBPycbSDTVWaMoG5Q7
R3M5OwGCukGpIBLir9d47VcT7LO4fwHUib51ezCgXwXX+d1xtrIlhufzviuknlCBcUd8BKQRawSo
+CltOJ7OmOj6otqj48i9pJZCquECwXHi5kgfzzHyRgop/z+ytLApz1e4uwRqiAFqJjTuvFHSOXuu
1vxomvTmlBD33WqVIjsJ2PURVMX9GfhHXuWWGJqTMmbL93eH26bXebKtQJ5X/EPXw43qx9VpS13T
R+iXElLwADS2p6OXZSFbBtU4JxdH0NOm7rAV7OV4atpeDrwfJJbBTZK6EWsfqD35SmNFPeOffvpP
Ana8HyUQjSf6yX4Ji4/Ub/gptlEt7J0Gw8OIX75yopIWi2iDZ7lb45nwDgfzCekEhBZcCwElQ3lL
A7+rs086I9riYsBgpFW24avUvn2hboOGNG4d6QBmUmHG9vYBE107QenN2h5ferXGQwT5WRXvs1Nx
PhGig2a+2xFNWVGzyqlaABtcenBN6EVbJhBprePsIg8x0mcLyYab1Kv1xbVPQKqM650mst4WwcKY
AR4q64yQuVrhOdXy/5EsiLsWuGEXL9tDr9L84utdGNDLRCejHrb8WZIX8V2tjQjK09L7DwMDI844
fX0BZvZfCsjZysePdtSq7EsqqkY8yN+ZqlTlDX6KHZFLdoiwD+mTzswVNg3o1ru5bVaGo4SbxRf/
8yq1EF80sU8Dv4GyIEwwtYy9oUCHwJYtObpYMttkCQShCr/xZbv7S1m1SuxPlE5LwBKDqkS2uhjZ
C7GbDKWdcGnrzRRecsKDRNCqWYVq8GnTsQzheYbUlsHSxQ52ObS7eNC7O34oQj0kca53du8SPVlU
wtWuM2woIpfbq/c6F1q4R9JvYOIGqToFfjmQgyiqT30Svns4zHzctfAN11A2rlBacWBqa+TcAkUE
1USvnZSwqb++H2+8PKSpfCxZKu8qR0jj/r3dSc2bftMNlQYXrwLLHUVMVoxIsZALMCmvQ+656KrE
o6pR8kNEGXa2i8Ur44KlUgey5JrYHOFynVFEIdfaLGufOqc7uRZ/DLytaX9i3V7r7HtvMzYCo1Zs
kP6tVAH6WO4Zh0Iqywq/aa2DVmYGTj6OkyqTFKmDzVyV2s4ZVEaQzGWyC/m7e8ih+n471s2QGuds
S/HleCJznCeIxGwFa+SRCwsElOvYRPJ/jA7GnuN75iyPeB8tKS4kx+N5HCsRy+OD++F72eBNTs3Y
7Pu4OQvXGX0eotixox2HEPtGQbqutSBE5zmTt1MvGb+yKNclseqUCVA/j71Im3F6+J0DKRsASvl6
1OhZXHBszotkvLqfQVRYzZdFr9Ji9V8IOp9HPig/JB6Vu6neNXNe/bTvH4wWXoygl6GhbbjSwhk1
N845F1kEyVkC59daGDUv7uKPRMIHw4UWZNB0FYA+Md9WyteDCYNcfjqrg/0BKucRpIhqPG+Z0m0t
s6nkLVwWQNiRcq3PS28TOG3xo+6mhgo9QsGb5dwsGXlcmbfUVVfJWkQ8+pdceyjYMq41YgYd9S+5
0Btv/Bkp5sPppwl9RTemm7oYI/Et76K+zajsKrlx6GmAv2Q4eRnyKEkYXSEovbJ2MZ2U5EY2Il4R
zeEn21jtIraPqx9cwERjKM7hBUxBjzMU9qfo7/vDYE8MaL+4O07p56bHtNXbZStB3KtI8o1a5deC
ZvfrJm4xsv4RaJ2yEFEfuOUFxE6dFWfrzovYkEhnMgbQTbMbowP6/4hcwMaE4l3DKLoM2zoYv+x3
zHf+irBd/4bLFI1yclfZHaPgqaLf7xXGZKYGyycpm5gi0WNuxqUhuyMzKWVBpvhCr48aD+AMBHye
5OKoQIgBqEZwBAWM5RKQ1VB6OztlH4LALwmN68UJMWxRC49Kw7vbpkhpHoMX3gGWftug2mi+mRzB
LclRtdio+249X873HoMWbjIeJz8qEvtctLE5nYzRwLaZawPgCmQvi8rDHSdhaJgqMBsLj7ewrLjw
rSroHukAwr0MBCrYRY+J5T+YTrcgVSF56rxSJPKETt8dZM3udnU48qx606FoZ1jHrxLDeTGmSeG8
cbYwP+EjWV8UJ78G/q5Pji5w7zc5aWMNGoO/KOfO3NuyWfPd3TGdrQ8ZCy5XTFrRRp9B6BarDun+
rAtNRM0/rFWHQsfy0i9znryn+yPSUMG3aKp9TRxX8cauF6a7E/CV0sLPpNg1wqPhNUeGC1JegKPr
ERiN89L3nFTvTPvuemmJDV9pGJeE12b4Rm6kxAzXD66HkmJ5PPfvK172/Ty9YjaBWllleC6P9+HY
+vPTBrCOyMrkCAzR8ufEhNho5g5liAkWeP6tq1vvdwDrAu670qpzXdnJFMW7aQYphf+9rKaO5gDO
/6JffEFGwNonc6dCz6jOXNfSvg12GzlCxsGrlg5AkFzkOEpDAAJ7lUniSQ1nu0FZWQOgXzi5uHpf
0+NmVcpJavLoNVD27vSyI1IrEMidT+GIbVCJPd1z1nAFDn/IOG0iS+DTmbNYRC16b2O+IBCfrNcv
Nonjq6FZoxbLpcGEtxoDn7QNHs1kGcYhxICAsLR1HBE5+42u0e7PYa9dFdcbqZ11nWBifl4CfDif
Rjg3zj9jI0evyzK7hAD0gkntaAPCL1KF2b42VH64teXwViMFGu4sjP6/EXYsHJgfTUZtm7eMpyFa
1oLSh4WeTEBviP5ACGbWBaU4x8/pKv4xjvHA26eOIQ1WYIZc31Xu51VQmoJn6Gt7LRKiuQlycwrl
w+90Y7TQ8hk5CQS2ZsKhNC7/VZFaGWdTUmtiQy7uAOD3gPSLGChLwpJh/PiN32CpwWak5YfHt5JX
X+UpvGN/G5Dfh6Rq9TE1v7eb5yAaWB0uKI2YGt7PIEpViRQ7SaaufGuEJwv9MwojOef2w/DcbYDm
DZ/FSsp/a4J298KCWaHq2jQMu9xdtTuCW1ZPK+Vq1i6LrfwpgmXmsDLLPZKLNlYPA9v1km4KNE5v
Vz0cT0VOf0QcRoO6gkrPL8J8Yh5r85bKKejOucps7bVsMEw/l8Ym4STt65e5rGbpk+kUlvNXYcnb
6ldS4aqnKcfd9cdxS+irLuf0ZTXikXCccos9ew0pRcVHug1mz7sriDOdLS+EexGHPu2hg0CHgU7Q
wR7cfaqV/+FU6k+2+mqnuRz4Hi6mgRCVrYmbzbt115AnRKobouE6dC8r6J0XUfWc2A2Wvayp2ZGM
D3AySwPFzMql0nwKRuGTQZZIbJW1xnCl3RSHhw6JTg9/lPdL+N7miLsxPP5IbwRjr5Ap98LGNgK8
xuiM7Ct6B/hkemuT9CnRzCxmkzuG5c70+EvEBqia2Ce13OgCQTWJwnegzA5sznahe2f5A3ZZsjMB
nrQJT4TUikQotU2PTbzT7/3ZQo0LNhj3v0QKoZXk38/+yoZ0PHIOmee+MYXdjET49DQ7UcuUtUpj
YNfTPqBfxZtwyrvdHAe2XgLdc+7HTba2NR+Aut5W9Y1dDH1KIbbehZ6Ij3Sk+7407ZrrZO3Xxz55
dAjILAwilccDPJatAF/4iz6eIJRtTVhRnVOjyhE3mitC/1kHVM7nFV5w2+7EKxUrZSR7IkgLnIJf
Ngip4rSLyHrlSqWGtCYm/WykfYUQzr9erIqB8BbVBeWpyKUi2fysXXKu1c00Bz6qzvn1l9t6nrZ/
wYuk5Y3DPSORDITcF/ewXGqPaGzfomMHnwrfrjYb7qihHtKiVkmZxsCr6JGq+y/DN4hwabkqJYEa
a+owRjZLvB/fWRgSmamxTSt62b+zOrewn5jGdft4kacjVUb7iIfJP1rcWB8g02RpVdc5zTQBr5l8
RkPx87M6CxOaxICk5/Jd2KesIuOUkBlukcLEvkDlfdlO4h0Qlb7OxsVI3fZkUyIP1clmQQq/4+17
MsjyscDT2oJc+1gsjzJQtdh9LWf94isTFYyQn85r9sLpfnr2050wKDegq9q+aKNAgwzn10gy82TC
I74dEGfLZJ8rA3dQAJZ/5Z7Z6jMN8dj0Tv9Do5BKduzeF4t7XVLOiqddbhLYGD+m1VvMwoDIGzDk
hJUQPt1cPkhPNb6mFJXcybHyBXG6F8ppvzIZra0kJQMjqm3xunwjTxW/vO8B63WNmKOwu4h7bmb6
aGkHi73LFuHIn8HQyEXP9LDIvoKKirA6MhUsEe3UdDzvDhHbzeeW6kqAWuZYZ7xkv389uaO4tdBH
BdJFS2Rx3Ar6lvZj1mMAY/ni+3wRKj/OcdwEFSOMkzOiZef4/IIZnKp/Q3n36MfQ0TQT20Bqt7a0
qD63HKKJGH6rFqnRK/5xscpknvfWmNRXv2KUDf2ma6VegRhc6w8QwE7q0PmLrXVqzkNGmsFganOu
bgTj0RQtkRbgfOCyVbIMcacilFs7lAFFf+R+i+e/K/1+9LUtyYgwIJuVzotv6L7czULm068Cu6zY
ryeCEb/SRmQqE3dcDqg+fq860pDTzo6VsAjKOVbzabkWrjaAAvWZDfYgx9xfT+TqpfEiX3PNTKgB
roMKi1l3ZnnlvOHEqca4V37vio64ZW+9anMVUiIF9b9r2c79HF+x1OxLYxkKtqW4n6yERtR4PfDh
HXu/kXk5RB0JERY2UBfFkuNQVrBnGn0BAo9AU1lXQajRATj8pcChxXB3VzVpIuFyk8/y/oOAoUcm
GRupg5gyTWREDkaUE3TkEwKrSvTGT6osROkXypQbMGHJJQWVQfnJcJpmF33F9wfBI6XGUWl9skfI
T+0ZE9kkUsMgQLAFhZBNSKLirU3r1+bk+AWZA9xQJzYEp6Rl7+LcM7zqtZbqbOwLsz/xjCWQFD1O
T+mYeleJXNU4mi3YBItUWUO2dreU7izmZ6JMoEFHH7BfiwPQlSJrIjOKYx0bb42xDJ0Ey1a9hTFe
WoRIvon9Ofj4AoakIuuQ2o+0rQCeSVTNQ7giUjiSoeFeuWRLA7QW+tpbtzEvvjmwoyvjRkycUIul
dupwfi6QCaDeb/qNT6ieCO+zZwEGo8mWs2i/2x86qvjA9JNMrvOgYolQkrCNXuPuTOt5be/m9Zhw
ywpeSjm2jNRp6+1zt5tTXr3q5DGroqPrg/9DIx1NOKygCGUGSdzxgzeJiDW96Y7pHf1NlYapJwz8
chj24llzb0pIeSUUSjaa2/po33q4+EVF/2K+nGQhhQvFoTaTrmvhxxUShyV+GmEu7GDMtNmtSja2
75I4xWZk/SdpetahFbTJCtejn1AGsmEbgg4oe8ca9rHAnOdt+INcVxANsJiYWJX7EDl17TG/S2rW
DewuuOr3P5WLVm0zAEOiCZpT+Je+x/cnB/qOwoqqW1pYEGb2OCrZcz76B8ec/TV799288QC46MWR
RHpngsLNQriKsEqMO6Kl5ml5+GF52ENGl41xPr3mk7T8Zmhh8AtK9K0KenqBd8OjwZuZnDAW0ByA
KtqjuTS9RVGXq/blJjxlUFSsxzggMEpbT5EBZsQKOheAvJXxOd2hRefhxj92bQn8n33bFgGRaQFn
0SqW+eS+iKyUzOH9BOzbfQjM65G9mO+lCwI3EXw5AxjekOUoQ9v3W3nRu1Onn7u8jvla1fDKMITR
eh3euToVNv/sL5pJSvz+l4uhHeeZueTxH/RuN8tu4cJ05XjfN0nW86ZUFhD5k/6kDGeDPFXu7gry
ax0l6I2K+ubHePA/ymkP8N2jMQDY97c42XD7/8Celcqxl36L4cy+740zOUlmJ/VvIhLeCncCEksy
16UWHbJjOtlEgQf8808XWKbT07y08qk6CmjwQn+tycsJSuwsvcpE5+6U7zMkj4SD2mM5Fs1/uXbt
p2zNg3pVY+RkAeWvA4dJjk+afPw5u1Wk9lyHzlrYOZva4B5rJW95AOG9bYCNG5Avm1Y9s544xpXw
c5cvAveZfAAxrYVKNN63lfuRzRzdblLGfW6A3gV/3dL1BXKa2OdorvMU/WNhHDTQhF0sGjnviGvE
YaUP3oZyxDejBknqWPT4F9t5OzggObWfc1FkoB+CyKSZENMJJ+CLicMVImGoepGGbGdXLQvNLf0l
2hdSkpzEyBdBvHdA3rgAD2vqAvz4/QDnBR9/woh55IZHWS/RSpaMr4TxT/ozjK6vjpKPLhLTE4bW
pygWlrJegeHavYmlx5iHAGsdneMST1UN9Z539/nXIt4+ub9Mk+XMybWmXcFQubJL7GmnwpLU9u82
AAsysnHBS/BJxL22jle/xie4p1qUmgNPCly9gK7Za5/WwD038S+aOQ1UKiC6yG0IveefKxgQ4W7v
Jgza4XH3LaBOe13mGuU8SY2KpfsARYmq70Y+Z0agmg1Fbjpf7Uo/GOalfeDr74WxgOH0QwiVTvSG
7++/dnqBXkyMCqWSLenKSmvqWnJA4BoO20wrsm0XYg3JudS2EyHKyCMkBV6ghnssrkXFM0Hz6KvU
cJawd5IeeBWapfOkap8Bqjdm0NGj9FZUZhNnOwnhfENQM7zW3574ECen6ebgdFS/DN3K2MEK639A
nyYoXKpcuzLE6qLz1W1mUu34sYoLpgpH6KDrnI3tgbXYusv7Yc6uoAlCAI+K23kUhKIiz9XZY9RX
v/dpgPsdtyMMEHLA1vcU8gWBODlJOrR6TDPJ3r1fWGNvzYCUtVMVtGLU1QQfo2SkUCgq5XqGtMJ5
XPiMlz9y2hcyDuiLB2Xwlx8XotYXjpXRJobfGAMUQTLrCUN9urt7c2vzR+UylZBdAgW3gUHksquI
6eiJI5XZZhKM7Mh5f0ZpmnSBxFPg0CT5LLjscsLFEXHx+GnrLaEO54aZWsFq3B5UUXwH+n2Tbsyo
PdVjJDW/uPB5JQxZ/du5oX0My545jyacn3xNVa0CtAn7yEjezMp8ky9rNXRvS3OxPr9VbWyyTBUW
Wa5rqI8rzBVcJrVlBOpFc1FJ+5i6j+YtHvoN0syr3E6hEG3+4rjNdWyPBAxQm60LWCRncuzZcnnz
u4qJIvDe4usSvEjDBd0D79ydiRKx94XLQbdQUIS0Knirj8Y64CC7jskYdQQC03ktWKaSZuOC/9Kf
q4j1etR33su1/6riAzVgOPPmIJ9PrctNNo4SXMIXrl5ac+5iwpR8oeQx8bh/cXhDsApNqv4gyPt4
DMdPENWt2zbpaodUjTkSQ/y5n+zG6rk6UORuK+9ea12j7PS5HoFGVDHDyoFufVKMQFj63+2bmwes
B5JC3SopJrDpmEpyz2+ZQPzccuVoiDnyyKlUFJrRmWUfBtYFh3aqSIyn0sAhh/+TCrP36KLm4LS2
4hgJvyUl24IA+dx6/INJ0jFX+RllMancLETcW/GTC9e/8i4oKH9uKVX3w2IMaZ0ikEkQAdn8/8Iv
deFRi/R0Fv4DiLqkSVUjWqv7gmLUSDwUhCKY81r9d+hsSo6hWNP7rmBqiEJGiJ8FWYFwP7zduJmh
ygsWJOH/gL9kyEmKfzM3IN/g8Iuqj49d8Zg3rV4YdADuIoGOYrrcJ3h4uCh8u7dkeB7XLkHWuYwh
KNQ8qWvdC2RELm71jgdk3TRviY6xWK4VaEo0xDYejidR9VBcJFQNAYZRipf4dTpEHVmQVM488rno
vA/jQHTpZptDkHvotDGTEtUQPZXvHdXut4eaCEJP9sZgruqWNdFqp9OLqsmbvNjZTm74BFceNpiS
PRLfQcPR4pHy44A+NjpmGtFGX+DmCRyQwgk15rA0SFmTAkyWAz6XI73phh3/Z7DQ53wgMJrvlJVy
C6kwB3eW67jZ0lOE47q4OqNFHqoQr/o5Y+YmBEMXdQEs7/FVxz/5rAnVqU4m0KmyZtYf6G4vY//V
Sp+9uXzf/uBq/QcWVsPIHXAkW4qJ2HzOUfvp3L0YqPEvA69hR3d2qHENjz8S5S5jRylF6v+pzK4j
gq4unsSYMkx+rCk8HdPlIssIOnJF+RQsIbY4hgO7wle7TNX+Cx8gbltvK/nKbMXmJZd30vKrhey5
w+TvMJUao0iOYRfrEZ1MawI/dFWypyIiOiP/VONq0lCtaLeqjZ+TVbM8kzneaoRwGFeEzwm04ed2
YWG+yxww8HYeXidiPRcQpUeriJYra5ZArnUZseuuoXoQm5NciNOZL6UnFTpEzk2lg3S1vlQ+nOIY
YD+xmMP5iS1VK2TQOYm/IJLduonMcLFRU+CrvWusNN13+fOVnw9IelFYMEKg6J7CEhqNapBstOea
8Idx12mxkQGtGrg0BcAgKnUqEHvXpEWfgwVDotbscePA70B2Dv57tcJr/gTY7NrxcUJctJlpS2Mn
cVPjCimu1yHF6tEQ7atUuwj/LdzAmDqN7p1UnTKKlGbEKQJSZOB4TCVM6UYshH+Tc7YwvT2mxTGW
FnRHCsqmbSWXVzGDEp/bXz4F1cy5HapL7ARfHJas6LnAoB6wMMQdga5KcVrGEJQ4W3VJIAhtpRoI
FN3ZVuEyhjOjU3LtVZd0Nwn716wsYXpH+qqOKZrk+sLDhOQTFxAv9+tUwmH9eIwlFPt4NatBiMfM
AT2a00lY8yDmuhYNVXi/kwteAERO201sYRgKhJiX4Gc6BU/tTkF9ID14rTxV0eHSMe1OJE/my0/8
3dLxZboHtVpLDjcoao6IuqPP+m8NXmt6VHN3xJZWJhe4dfBBBVnNjJrwGsRrv/ccukzjKfhZWBrI
6dQUwph4cyU2sLDHo/h6ex15BPIIBS/BfJq4oOS8BbRWN/G/WaN2l9fKivpKRrKXizILuawt5reP
AfGPrG0UZPGuEEiorw/l+HGlZ2yuBgmrpgWxWZ2wVh2HB9Mld6JIgVuVSLJwYWMVQviuKMFUdAyf
cuvivNEKrrEEkz8asU+lIkfz4zThUgPaivqSV0yTBTRW97WmTo+pUXbylKFoq2bfxEzhwoUK6S3M
79yV52q6P7WTEoW7wTM0asKczK59OSLAsMqTSNVBLpxeaSj8VbhQIEbUEaZ94pzbtG7nKusolSA9
dVkjH//tl8elIZNNFXl3T8anu1alEscpY2ttijF4AwcrFPEnl0dVAu+9ZMUgIB08sUaeRmf3wxnV
blEAJFCgpoJyjNVeLsPndR2UHkTX51/sjRNjAP+2fJkLfgau8sf//O4kOTTKKUK/fi01uijuPW+s
zIuVc82XQistjf4U8nwiMovb77HyHr6i3VhGKGuPt66GqRKY/besHhcjxfoXub1HZJ4C+f7fCpRr
g9sGmh6BVX69Lgdwz2C/9sh3041urWSjX+HtPfYpx51+WVHAJ9o8jZOp4WeNSl4wAS9oyzx2NKZI
ik9gBsz7FcdpPmXceCJc5Y191CnBsGsG08yde8kCMsX/RZJ4dE0Lat9MEm2RHo4dcTjSrVt3F4kI
zChXxxD2qNt7i38ldvWpnuam+T38vb3hiF7v7DkYTuSslwPNSZ8PyLOhGtc7hIn5YFzlq+NiXmxy
7ywYZ/57pGaf63m7PIxGthkVx4EvfctP57nVaHIizAsaeIMG1IQjbQmdmof8mh7UHT+R1/7RcwyY
VwRDByTYzKHJXxcaxfsIUwAfGkOuk9LutjviAR0rDRe3UuR825+w4bSRfwiW9s7Somnr/J4SiSO6
GoiYMlk7l0zuDb6tNmpr/pDuEpMbxyNdin713SW6xKHIhJCLotFpyd6nQ+zhtlEFpmsbZIA/TJSr
5mKTNZkubWmB7ne4MSsE1Hlfnih3NnhwOvFR3/Gy1nEtQiA5dRXUVAbKu86iHX3Jpos6PYP8Rhow
WffUurTeFOblEevHYrz9F5BQo6NeiZUH989KqapWpwZWDyCMV4bXNR2Om+zGqW2fgp/XG4Qs98qc
shJBNww30uqQDo2zuncJ8vnCln8QllRoOOp9EjBOEVXXsvVD0KZ6hsxa/0CYlWpMNwQCdgE5MxOe
54fy68kG4A5wSKXvVi9lspdpHlwQZ+YpdqiWkQL+1VCwV2B7ivo8VSOue/dJcCzmJAk+A/oUirpa
QKum7e1jnk/3S4YfV4MErfcXl45f4sFtjPT+T8e8EuoFWaV/flcVbJklBNizZYKQUP7BFumicExY
71W8dGw3k5yy4oSwdnF77+M4CWrnlQz01pGlsgBxoXtqC2sucXkwth5pY+CE5URQTLWItepmpJol
tWtP41SWSFZr//dRmjLYUwL6q05X3L+KmeNp3O8X5Ah49OxdiXj2QkNjKFWpgOUapYnyDP7mkCQo
fe8jpiaITw2WO+76Fm3pVZ4gl+C2QLZOLtH8zLg4KNVg3pbCoUJRErP27Ksv4t6rLVsFrpErFdrm
rDyRscN+8caCtQxkn+GwC8eRdsBAChU7fHXaKOtTbrN62JqRAKj3DxZrWKnUTGVe9QxKpWsKJIV8
Q6T7EWuGTnM3gniNqKf2kmZLFYWLe5bygD199UtmfSiZ6rQjTgDR5lA4E/W08XPD6QhU3OfKs7AR
05EClvJ5hi5FuSXa/IVv9wNlreZpP9fumFFLwaIZGOTAvw/BGO0SiUXpax1pZVyZsUiQXBouIYPA
GfVSpZ+KwK+c6Yw97F9VEHsgCgVMLUK6fw4SHEriEZh1ttmiOMgsRxUjOq3UFe4E6aZUN59fk7LI
4OJVAE8ccGWd/LXSs/cvBdEz26vIYjcvivMHRPxTmp/PyWs+Ygtt358EFHi/9EmGIpvW1BRElTH4
pZ7bYtOalp8+3eE9qgBNS096y0pVXif/bjK//4vqqQRJGphnS0PeoED+ynIPPLmyACf7JPxeJZfk
DoVCE7VaKpAhRl1EIeGOW8HG6+PTxzWJjMzQ3G012wVJJT82asu//hc0d90OCak5BhlTriZUIyEI
mDO1X4E6M6gxAS9cjWWIQfZa+wNRGzQHELu1cTr9gfdbfSbM1pSQtLBKzh3FsvHJIg9cvcj+A9ip
radwYuQrTTNIqwcmzyrmnksF3i33UbDzraLl9jdsA42YS4kK9XM845tpFJaXAhhc5E/GJCrkZYdF
z22Isa+CX1vAYYTa+bixjCvEpOIzmFAybbQN7P9RO+4vFhNsOHMDBe1LU8rsRiSoUuoGAmLTUGj6
NLAk1R6brNXCoFdVtcl71Irw9OkJUKY/ebfYPiQzTtkphT40d2mEjneb6lAgF+SyOsmMlGP4DhOj
VJzGI7TKRP1wyUapiFOvNdsioWO6lzcWw3NGt5EV6kfZlwKFwi24ZdnZT22XB3/61ugxta3iz14T
/YfSC4VSjTizUN4TtEq90dCUvxmRV/DgnKJFNFxqcI6N1RHmq8T3u9WI0elWmLljOSZ5GJ++d54s
aiIpZeeKRcaEM5TwrqqJFrUee9w3PvDHe6TgxXLvusH78eBbdk4R5sBfg76Yi+yMomABJjXiRvPS
IZBlcDpNXvkP4izNQTgXFirzEkNPKIaDPUp09oytJ1AbGOm79VwGgB45H9JvabRY3L52mF27Kvb5
sDK8bl1b2SgDPW818qB7GlFgzSL12lFuq4PTwLN+D7aEYce1+J5/7xahAs926m3KPXAFYjt9k3ic
6c1AbQ0lqxLGnBojo6Nm2OLWAe9TMmOrXtkS6ldWQgohF8g3B/g0eWrElw6iLq8XvHbHcI3q6DnH
1RIMplB7NPhjGYIKNpfgpKBiu/Og3eqOqH8NJo1cabTS5wKs/xpwCMGxNmVPNdZFShg1hNBmUyJ5
4+th4wI0ozN/JFYSiv/KCyFx9Ht8VtKSqPLe8H4onr64HvW0kI2wijCNWdidDSTSCGDGNbdG9Rje
a7YvifHS1l1sA4TauGE11oJtVnzFuSWl36eMSyIyudSj6LLi5Dgy1Vi6iq6V3+Ovv1N5Dh+ik7lV
eeElNVXKgxWUDyU/wXtYOwKdf/HySvrrlCUvWU1prbmGzfEf7wpSMn/bhl8giEL4zlXKYAIb1AKq
7iWEzpQSI4kQOD6S//VH5oLJGfL3q1ZCL3jTy5hMu6LuV9Kbz3AHdZ2/kA2VRh1O3sP70MM3Q29d
EMxvXPBT1yCaMVBt2R/DeLf3q/sJDx5wdno7c4t/5KPXGO/LEtWFn6Q3LwAUaDP+Ejd076WAEywH
OfM/4iyDShXKBPDSQBa1BxvtkhECeYBeU6MWq5drTohzidI3TLkgsOK7fGGTqPW/lIDEU4BdQIEY
OxCK9/vM0eZEggUkSR9nkn3Omql3TtMx+mwCAU3hDEpv+p+r0fz5Vv7kYHGS/fyL+MLJF2PfDlug
s6ITk2tZVyTlFJS9uB8GiMuTgNamRcpq6w9BHf9s7B7Xjc4uNX7XQnyDd2cdBsQf0YTe90zpljrq
EC152VStfiAqJafzyU48rI+2s2C+tj1c1DsnEpG0EiauHVJvBM2Oh88VG1ZwhXlWZwxF/O2Ok9OW
sOlUHwpida1xfqExfs7jz+ckWtlMGtns8dKrdf3ePWtziTHa3PwTZwLCm+PKPmxT93ckBRPo3XDB
BbGQdy6pN5aHfpKFwpmXYL7XNHLvZ/XsjeDi3/IwdM1bsFzmJHpgxgDmkzJR4P8WP80lqltls6J+
ZC+C6SxjI3Db2uMMDWL5v35KBTmVxHnfBKPTap7GGZpOqf/7nmxPDeqBo6IIUjwJIqrJEYRGBmJS
HU05PGSr6sv6mAzpjo+PQsJLgE35fxit8IianWsMg9mzWPQsdWVwieFq6r9UagW6ZSYYdYEKKtAZ
YyCmQlJruV3BzxIWQnP8aE/33ltax1Y0a5fFNbsbUfbuRGa+wfaahh2P03yBHOX8r9KlMkmrpxyr
HAGtga10xpxgVxX+P/Om3g2wYGNj1meQZVdNy36cKI7g2fSNYXsrHTG3ue7a7K0NsfOOEriJdiHu
2gYsGXLEIUGW7DV2EqzYuBa9FTUteeWYlaDTdsidqMXdO1JOQcHLDpZJ45DPTg7dExU/b8T61Ucr
36bWerkytuES5bv57ogDyY7xfX5ks9g8QAqXTZvQs1zSLAkOvp/cDYLkrKBDi3NN6iiioGp7olXz
T1zA1O6xGrziTYtFjjXIprbt4mMQdvylgyF8tzADUBC7vg4DE9kLt6WobTCHBO98OepydbXUfzoG
ims3IU2TUgDD5Lf9N+46UZkO3gtqmmgdmK7a/cDFI/a+DeEbex7RySfKjt3S650UHxcRoUmm3ZOW
hyJ7YhVOm0XOAL6Wtu051Mlb0cy+c+wNNXz9aIhVGpocGsbNJrIOUlS/9/0uzpxgfWaN6REqOzOP
JCWAXNI8nHJWmgpHz1G5PsDmvyCelSOIRkXpG2AtN17PI33igugYO6pzHhuI26AmBnsDm3RPHbF+
MicKwUjsPt+NNV3B2ijSvguR91op0n66jokwBpduMf90I6WFPg4QVLDqNwIX0PWWPuf2uX6gAWKc
STcFlvy20xlDzEYlC4t6fwjmcSpSwhTPg0mD7IduJioQC0rIhtUmVmMuG6X/CTDZpUQdfPXyldj1
56A2fLTKyIHFrT5FBcJ7k+Sq2CR6zULXSesYPgxe4pP/zG70VVmbXsNdXWsESOyn2gGJhk0ljpcb
vXvRzq8/3ZZN7c8tCOaXKfIy3+BvhuVLvTucrQMjuTy6Te3FtgddMA392E88oyhm/soHwBcJHXbK
SFGUk+iEfohyX86W1920I8A8s0V5FrLDogQps21BN5JB2z637oTZBLWNw4AY61qzHXJUCF5JW5JV
NCZEIIIMcwPAj50nDgpDmc/T/LCPriSq35ekEXFvF0eHSP8oD+iyJtAbZ5ajy7kLdoDv0ifQGXbX
AzNnhRy8Ox0QigVKKqmCcbVHmDJHPpkKPkuOs6GqGHG+k+Bp+x/6BzlSJoUvbZA+eZJcl4avS90p
ppBA+C6AfwhLqrTsB8hWuvsddKqv+K0E6WWyIAAu3vgIX3XYtHL7cWu6rFFhnOQWY+qpK7sZNaaA
jx82/PQmFU39ZbKeQj7uL2HVFEJ1OHXiOKNH9yWZpEtun3mib/2oR+ZtjXCbo2a3qSMX86R7Gg1T
Z0NglPczuoDhepwg+gm4WnnD5r5f9gJ1tSyKLQQuU6DMp/y/E5u8q7TyOJkwX3aXOixTrdFNv6pO
KzhqG/MWOvID4CpvdEXjhHkuX4NR9KQQjJ967wEpc37ITKDut/DE06pSTlaAm2qnF1mmLWteal/+
dg05LczCVFFXV2zP/dueb9Vq6ig++r1kbMcKe2wgTz6gO2xZfdKGodXL2KeL4WqwFo47sDrEcSV6
kjNMAqzn3/afrsI3MOLgXkJ0HxCDr9XpFiuLwafH6bVlLEZH4N2amEQBqUUpcC2L4PWKFZHkg5Bg
chCYoW9BA0+DR/f4nvMC/OqZTamtdVLHZniMZInu7fpCmNx/vQ5UPfM8FcDeYbwTxv1hxpwQqJh3
oBxgoDkXeTN1ENb0OB/VpyNyMkuFzkBPUEmsLXyCVSQfoLefqIbD7ktCNVhMjtQb8VROZhKtjnOA
vME1AyI21Jn4aUgNMTd/1JRAtLhBdoZNwAxZmPKN82wgVnKPaMTIq3Baj1vRig/z9f/YWPy3khOo
RX46SY0C62xWZYkUo1fpucf8wKRh4cLuAOzK5d5cGPVZ1ISetPleBj81GeYdjuVDTpbbQr6UXBAC
9oOxGaYvHX4lVFq9mLdg2zFsaXJ6WKdSPyqzaactA1nw1FWQBnigarEJoP67smsNQOjNsdv+8dU7
Go0jeGkXZhaPDyb/itPNcuehkIa3X2UHGLXr7PGNoH+0rHSgp4xOA9uwdLOUtxo4nSpLPE/MojPi
IonesaW58ngPWFcxTuTItp5WeVkIeTsFryknR1IjGeh611IohIy6UM+A+vIWXFzIGOkxJoWA4TUV
Q0mIyZXOyR1eSz8D+BoUbT+SV8SPrcDTRVOwfKP8JuAXEiOvg80sOKbKEUPQ+BAJhoMg2JGjTqPe
2oRiS0lOj2QhWJfO8ahpidZABx7aa7joyd90ooxhnM1EfcFLrJBP8FS48xqUAwlk+PwOKs3JgiIW
yOV0filJCFsS6krMD5NJCtz2xNqNssNcZiAl9oCuNgFxAnI2m5cxX7PgMjd8acEcOl0EAY4rHush
OCm0VgClz0QWWdI+E2kntDwJYmArerlJBoLwrma1oVheZJUFXS4niyNo4/yh4pnM6BnOtWbMELRP
sAvoxkimYnUQOpRwF2ja94GlIEWI6WclXrtnrBYvUqSEHEVXjf8h9xHQDB247y4xqRGGIwXV5v/F
+489xyBObFAxrTGlDZU6TB6uha83SgDsWydRzrtKaFqOLbXwWuGFUoN/V1J6nQNo6KkdwtjoWqHh
YW00HCHYNDYje1CesJEiCJkHuPPm+7ZK9QzN87BSRKcyJ6FTkQ7HSBqQ/sJvzLC1FIiXW20KfATf
a4sFOPTSXpptG8IUw1sX26SYZFEIFhZk6N9KzSa7pkku4G0rqjm34oiL04SSDMiFZLVZnlcSXV4G
R7NtkRR01TeFR+VGBqcc3zueMb13O0ezwC1fiUxoM2ouGjaqtrfzVOctGPydPx/apem9q4TXaOjT
KX/l7N3Goowm/zh0GMBsRqH4q4f/i47bS0tStJgSMcbWUWukBtt4YKHoJC3DwBjKr2DeFkF8ms14
IBQt1t0tZyN03M3Xxhkz9OO/aKCxkpwcbecsfZF9CLQ64cWVQAGmftCCmikTmAXTj1Jk1T4uQzvO
Odx89JMjDkyPck/ejUCGzAahLnVOiCKiM+FaCI2RlKiyM6g33e84qs4iJtYMXOM9BiH0gU+D2p39
NkvIrLKRBecuoHifnW8Ij8SB/ChEtZpF+9DYIEpJJLaarbesGPdAKtEwaeiIHJyqIcQA9Bta+SvX
UDLSo4DskxQNNRoILyxr/qfSgtrNavW0za2B74OLHwKCZNVRSKH0/OCyKeLyOj0lnggLnb3ws/A0
oXy9YD1GVKrhl3mQBVuTuEbvo4tOkAITFnttUI6LtKv414/Vyw8b0E6nC5SAeDQbjIgmZzGeNX9p
XDrVySp6SBxw43b4IHnYP1f7VGy0a510zKtj+9A1gqcpVIWDaU6TiPuNOJbAnLCMbNUUW71UJLtV
IUoq9E4eLNshrlTo3BK5hLw56AjcY01nbnfWnCl3pKnMVJ4bWtsIVfhu0H9u4By4TYxEaPEnQ4gX
hnrepKF2LkB3djXFPn3B8v/VDR43BuzGETmSYJSKBQTlNn32sTx36qFqbV7Q3z2/rDNqyFE19sJm
SCw1Ipan+1HFdelDYUXUg9vzKl7m4ifQY4jwSaGhYmZPqrYMIVpnldgcV/BGGuoKeYMFFtWuXsvE
rry1BFBZV7Wp/7D10Z0uUJWFUrCwrTqvoKnwEkKfj8CnqjxyIJ7eLnlZNCOFUEE9KkHnKUHI1DZq
3slFDBVrHX2WmZETt59x6uyek1Vng/jTtekOPgUtDuyw4oFuC9U0z8vUTYaHQzr/vrtfI1ohGtfc
v+LdTZwOjRkILRG8ml2oY8GxiVQLPp1I32Ejl+Lm6q3KgjlERSUjyQJxd+FqG16Bel4cK/29Q4DG
wapSA7XHjtJbO3uZijdifLkp7B2TlGYr7yuknDKAvZBII1Px6SDDHIEfZLrfji+9uMrCzw7rqufa
BodpRvMzDgJ7BAFNmskJ1MctLfKqwDR0h2qo0EWmucmR8K2rUsAXqXrqpWrsoRkv0oGzetiIkTd7
ApuQ8c55HHojJ7HxWZfAzp0uiq8v2sRFoihjyPxKBZZOtWZPJ1sJP1AxeN5Rx/TtWT99OczrDNnp
6OVKiU+pky8nRLk/KMcPdwZa2Wjpa8ziAPta6yspZgKr6z0Axsg8oNxhUeZum/VVKef/yZcjRcw1
/0E9zZKHrm667+9lI7qxghQ3R5Pq74tmgjXpUg2hhM/0ZyIXxRWEHW8yvH7Q4HYAUr098TPLZ+F8
prgmv17uHJWcHJ7rk40RCX7inlPVShRCwV6LtDKRcmB845qgy3vI3ch0j+v/CajfDup5KsroCdEB
eObt17avlgJmrDH1ZRZy/A2Nd2a0GatNsODboY3uD2MTT+xp8IU12/k39185+5ae+bBmP4JdT0DP
EXkOye7U7Aigz5qNbTge4SqGaRVl+3HXKSk4T7DkVxUhHLORKHpycPx85yMtTR/o9Lp5v2TaAviZ
4xDnn5KCBxu7Gcs6kKRoEpqxfsJNHYz7YOlEssuZxeLfDpLvUdaCUVHsfFAjpG4y4E/jpvwjfOr9
DI2FmEagRFxq6gWMK85rt1aCqDq6IRLh+4arUcGjQlsGqjhBd5erdQDdiP0RbMS9SKLPCtWlz1Ty
8edlrb81kHXadNh58EmYtDjf8C/dqPJkND8AS4XsfBwobjsJy+JbAMv4WV8z8wE2QVtrtcYzbWAp
6ftAmjV9t3Zcn59pwYAtp0B/mr80U2SnvxleUBO6rsL26PUlJoDyhOmIm5xvZbH/wpLWY7qlWz5Q
sFywOle4thsbHG90gdK1dJnd5lLdpsuA0nsDRjZtDUBOlew8DzLXFXLk58ut9frgYLJUwKbi6AdK
wK2ctBKkY66CoyLFn9U2uONgermDzrIpNtSuUvmroACiHsUjFwLYT5qbZyEp2NCPDOxcriC9JDBc
PQDGTKpgwTmwRdswqmRUL5tjSpq/THy1v+jk3Oyab8uG+5MBeRJt8CMdtgCTkf9/N7sSJ5yno0SJ
rpHwng8J5ibTlZIW+3NdF/I33Prv6YoGBaiZUWz0lXuMxBeSCEQ2PyE8dJpxBdZYm4gPKDXSAO9M
u/itqSy1s0rRzwB0+jhT6FiKIO8iKCOoQqVMTFBhZ0Pspp6/ljm15nkntJmgD9Iv3TRxxJHw8zvn
0wYPe02kzCfgvIkfsmKl3dMomcH/D37ZGZA2vZmhJXleP0fz+M6hj34/4awd+pPkvD3IeXJd8Io1
ygBy31kZzf3o3wNxSyWuHcgcw3hb8TzEEAJwbKqUOA7E9YAcwLoRc/bc93YSQfZMdRNHJud3GCy7
ds5c4xyTeffMAD36pozAtEyFz4MtMtIzAkp0NfXHyKVVOBbaLrmyoKy42VWYkK3cPA+VY/5yFJyg
A7W9hPWsOOr30pSnKwN6nPvAgdSNRkeA+yKPOETwXbYY9ofdISC/uSH/934nNYgDOzaQxgusCLiY
lOvIxNeyKcJF9Wo9K7NriomYCs+e4cCdwYP120EJH1hN67Xcxe8X7NvMTlp5jfinJkwrUL+1LiUf
LmKdWrGIEWO6CVUL9FwzqbcsA9Y0ALXHIaRgKzDHg5i9rN85LvRk/2X0LHRo+Oyukr2Jk9jjJBrn
A//0xg/56hWrfDzNmJSIDZwsnSxyt9/sh6+LEW+WNuqETLi7+6j/QnLZrTJkS3wNsWdqqt8L6pk5
BGVHqXya+SU8jFS92pYzwZL2kgDX4Akksssmc3VCKD0NuFGK/Gb76GwLtAkiNr5L19/7UI3lQFDZ
AxHZQ6XqRDgGDgcW20cMcwdVn0tboc6ib5eRWdlo+Qw+Ig4b8Pk0K2mbs6misjgGqNsnQWqYjvuL
CbjTkV2yrf94R235CA0zrdkDJq3t3+KS4o/4euFBZJK+BvCBgHdKZPf9Af96cwdTzZpqSyQLdUG0
qLhpNQVzNeE71lIOw/t+RnC1jFTEZ3qaN3colsZuMxeFKQKVp2jjdRE5mxpt0VTygrI1Fag/PGUg
TD90WIuD+2zzkuh7hdbt4OehpAftQqPcTRrBpHqPH6hVxyFewR92JkukCcSEMwIYRPpOcRFBS8r1
xVgyDgDffCEZvgoxOSdK17NbOr99myyjzaUt9/l9mbqNlcgrS5Yl9CoWAlX8+62WXN/SJVCUTbyc
jHU3LzQqSLY3luit/6slPFQjFekxNegR3FqfxT3NMLeYz6qbUcmr9v2g3HKesDpFlyZCb5NFY0H6
LYFepP2WEOlNHIqUwjLeHs6krmnXasOq5p4Yf/ngV+whfwXcoyXXt21XNOMUVnaa19ruswwYQR8m
h2OgrTPdcdOumwE2BnC8zfzKCXXIHM797m/07+bpufkkdly7iPGSmtRaiHiFd2mrK/um6nQsFcZO
o6rHisrlJsPqYHqTUBeYQGncDnM+TudPuQ1oZGL1QUucWh3jmevVNBKr+3jWV3ehDoNhRhflJwoY
TdJx53/VCL/8YyGl2CXBN0BGtOIIA0WB+ORzh9E3+OqfCODzALPqUMz+wz/q2L2qKzMj1tbfh6BD
a0Lij1tWO26chRkfqVCS23j79eI085J4l6CZcec3ydn3RSoDdnfy3+ixmwtNNXU0vTdqUPkEImhE
htBVwU4sVQwwMKteX6Muy7/2+PymjpXZRAGlmY+DWnBc/jhaFJN4L8iDj6S+GVZIYycD3Cdl9IHL
CJnafKbOoTYN5LWiKbgA8jqdnarG95WdyF1Z6gB0FibKlcYM1Tp3ro3bgODXkXrre2EatBZheqR6
/iktJQdQ3iHnU4045ANgbniyvroJlGvqexDyZy8LY4FQYr3NpC79Qo56vNruwHpoX3c7uV7N2rSh
miQSZ9xnFiXKxWxFDbsDD9DWZiHBf24f7IjdhP6iV44M1RBC9OBHC1tJHaR3DouBzIifnVQAIJAF
FBP1KZ7uUbeXlDrF6aulKVi5wi0EK2kUVAC+DEGxMRpKtNJi0C7M1Y7xp1aQVuRNBD2HPzxRDRN6
ZILmw46ltF0L7XXY9PY2LNlC5v8s+5wfnraxSSvoqP7/tmvHcBwnROnRZPb1HeRjdAPDb9asjA1j
+/I+cBv2bNhwx/zWyMc0yVtLOBwjS+pIZzfaM47nQzNhzZIRVyLReaYDpWtCboXlrFXb4i3lyyTS
Vym3WE2N/+pydFowwMypSx8laW7c1Peuy+yGD6RDb5xXyCNmoVTMDGqk/Uc1cammr6R0/G4PlA/Y
Eq8A8CQVUMNGL5s5XXrWHA7N4HQyzNGvLxjSoMDapawXqPjvvp9KghgJN/VeKQKHUOqNh0vtXN12
KKghVX3lVKSTedE+2tbV7VxQL14jbgYgdWns+/yYSG5VxBOsegLM6blLYMmMmWnFIJV8ncUQSwa/
sbltSxc9HoVT62ILPoNQ09zVb3Wn5gLBISiKP6/EIYrEUdiZcWGV+RxdSx2ljJjgqaLiOXHTKGPS
LbXCohWm94OPKHpaMpVkivOshGQwwQ6n/JoX8liS1d7YfP+Nno0XMNyG0iHluh1mHzIwq9w6/99+
g4AQNxfgBt+B/VKQFb4muTPEKrueWbG++LqRYdb8KpSee8BBkEVACThi1sfiESMq0JCjW28UW8Nj
/Ao3FCqBr45WeMTwlHI3beRjIvOOrRTNr6d99Ax1rffborRKjUaDqyDO3j2+Ec16uNdu4krmcfli
twQxl9MZeTQKrujY0me7pa/pGOgh3AjHvlhoZTMPXSCS4wveyL6wewYDtsZknwb+s5ibnkjA6T/5
vrR+gsZr03anbi0rkcVE6bkmDF5CFM23d21E9NEHv9pdKGUU38JJn6AWUN6UqLirI2q2V/RBOsdR
OyJ7EXMGnVYkLZh1/K7C4QzGWDuOOg1s87jf7ykJERGFbYkhcAvFVaAYPmT0G2EImXPcBnKR2aoP
g7Q3TuqnHygF0hR+v/JmwhzTDkaBD0RN3eZbGj9KrbQIx9mqCXkj1yyS2fS0ertsw/vkk665Gpi9
tu+UDubxaMzmMj3okPFcH2sjdVQOH0Z4y0ViTGpI3xFLruSUhDJBKO9RUOdr5dOiIh00nc+HvG1b
mzMsg1AHJ6CG/nodu1+Z0UXFOen3i9M0Qxcc3ig4J8DQObc5BMP0XSNEB7zpJdY2oD5ac5PMiJpM
NsVOhV2oZtX1JbRboUF98fefo48B4sjd1luWMEQp8QzCYxk3pu6uWEjX6woqfLMSgpEAoyKxX9ep
uifaQ8lSXGRHVLIZDJcH3/4aiWzKrwHElw8u2B5ZKskj4yT7h4NML+bgrvDdvpbt+FWXIjP18Y8M
KHIEDgT0ThssZgDJhIFLf/yB+oEZNFcPwstpx1U2d8FAKU0S654Dj/s1a/2Krg/9QaG3tS9W5T3e
1tk6Zo/ktu0sg47EjlsLhYUeGE9jUJFXdiPzxgItxwV7whEuqBzVQFQrdrIHd2GN0ZjHVscd49b5
LuBGpG8/ndJtEoYc+FinZhdw5tVysUUWwYEEwNb3LarFB0IIaGxDU89+oEBwtyRgnkVJSWXkI8pp
qIvucbEGCNWuYakwjVKEfU1YA3MqsTl3ciI0pcHz0OsiGAt8wxOf1nJ+eczazmK2miTOvVtFTa7C
NooT/mEsNh5uSMoo375nV1bIDSqaDugnmDEH7+ey6vg5AvApIlmbkBAmMvq9ZrK5t/nZx/ttBHdC
nwTd6XLHuuSGeZoIqhQyFplODqV1GiaSSXIBOBo9U4q2iuve7JU2NxpSJjkkQKGnmGvPWLBAX7JE
/uUgj4YOzhPQmUz/HiamwMHi22PEPs0VEN1juGUOR0ayfyqHmhaouc8T+1qQS/OVFA1r3wCX4tYA
fKC/HXg2fkBoKRSI5sY0CSXlShBlcCxDO8WqWp0seXC09rXhyWPWf3mjRY83TzrAFaRwc7YL+WZN
dl5R5uZk4EF4Tsma8ICtRyYfRxdt4Kyhj8/IhmETcJ4vpoXJTe8jH/uEiFYsr/AjvI6N0j6ZWiXL
CEKCIM+a89S/N5Lfn2QVixDTisgiX7fWH6j4vwyaMkVeRsY51P/S6C1f5r0nRgVQr8mA66uUphbV
fsAxqxWO+r3BX5EtmpvU7vaIjX8HV7s8dcpWVGizel5mLrcjY7LDcXuWHGoRgtd4x9sMT+pyh4kl
6JdI+/2DKEpV0CleoCe6SNFYOZ3X3tYmW7RZHxKnKQH60d9CoeLALw7C+tYUOvwyXVl8S8gPpAib
ISQ3mjmjLrO/bfJSOtYKo0cdLCPJckAx6jSApHRZY7wTFp/rpdzTXBfw4JdMnubKdTxvk6NQkQXn
u1B1LYW61V1vOQOJUy9mTfFJmEUWvL/ujpr847Kon4NLG6lUXtW3ONEiqVEVWzcnOVWrvZaZd08A
kVG3XlthBXgyNvZgBYNKdPa9bSlAEBOQa3vZJbX4TWrRKjA9eA2zCiZUqcEttHp1vT9/UNnK6NOI
81M7HPBxg2GN5D4/M3bPltSwqZ4x2mwsRgXAkUYxd6pzT5AKrYCWhS7CB1+9wOHrHvZiGKeg0giF
S+MEhJXpVMqjC5rEdGzLoEEHdZ8itnl7PMVo6O773IBf95feeDN8BLyRFdMJNIWKcJy2m/HcTmrl
AxqtLW1PipBOoK2+Ii8RR6FsM7Dn33W0Bu89HCYwzqZHdGBup2ixuJgKwnQSSdHCDryixmunYwn/
Ti0ysahhlTiMLIb2fRRqsZ7GgD55VKdi0NdCMpCxXyDWJDjPIjkcs5VI4eRQ+fi63UEXSEQBUSla
zxC1hSljYBtbi4XUhvuoxII90VJu+91f8hwcuxv7JuCeMell1vr2lzoi5YMQW64MPi5DONBAo+3t
14hYYMpaVe4iJao0BDOhbd55k8JNG+DGpidv17N+hw17fHe496WcWCKijYx8sYHaDvxPNlU6Z0o6
9Op//qBW4qfUuwGfHa6CH/e2pYUqltBgAftmvde+XUYbMm7JpbRVD2PGzjspJXYNKdQWu/Ph3OEH
qpkLpfdDfrBKVNZyeJUCLG3kMJ7iU9zoo7EM7ArhmwKZQxTa+owz0tC+9x9THGaUqmqHFiOzN7Jo
5jfgiB9oH+j+9fDyTDnRiflOlJY8Uct054xD/mwaSSm1BETzu89I6kUvmkcTWyE5EDEP3twXiBG2
443f+irpyjElPtYt8Edv2z2lHlBgXfrwrbYbg1VvgZXJB24/VRwq34crNZVSyegMYtB8bUYrvD0h
ZQ6ZJr+kHMbOrKr0a6YRaPBko1zKB662KkzYUito5TS29yri/uLtz8bN9bukDmpm3iigaAzkvozP
poQukDSaMgCr0EldHNiq0y4xb2tNXVdZvChZEV2tWceC9RZFA1UY2TOoGdYeMAVVZrOXtmOUj+vV
9WzLaCDl8ZwhV1k4nOdKLJqU1QgyeL1NvOjJA2KbJ1XYrN5IePtmPdCgFZcPn6dstXmLBC6/dyUM
+49azcbL9NtB0q4BSRwMmqWtZ0p4rUdxlREnZj4mHhY2M3pK66aWKbi/OPkR2rR9mjjyiPwfA6Qa
PbAs+TtGQueRs1XrFmKU1Sihl6+zV2MBI+R/XPz6D/6bWf7jB3CgpKeOikIpAFxx76pi/2AFYjFM
at1WLtApF25qfgzXDzag7hDStP2f7BknjO7WNxPHFpMVJo5R/nSWFzYH+5mhvQNmLBKpT1IwdTTV
mGJQxSCD8PMsCilQZFmA3hDtmJTrFGW90RymOvV8obpRhtXe3UeKir4+ye+22FEFeSy4nK6WryU+
xZoHBVUmwH90FFtL4Ah4Pw5EyTxf/kHEhnVIwbpFmwszesSi9UJlqjO+RKSNfiXSEsFL30wJuGSZ
gvBE4F/mS7NNbW7krwkUY8SiARSvcHdOUt/lcfs9xPlmhwxP0HjEG1rewDUMt8FPZHJYZt6tSnTQ
y87PpT7oEJ1RBRKbnd2BwTIWp9aa3dSbquwZvQPjeogdQR501zQLtlDVTFH6Sw7osMnxPsV4VBwb
fRqh9KFvMhUDDx6ARK+WIjRFzfBpu14EijjxRknQXLJv5eadtyh8q/7p2gXFbQg7mqX1kugI42rB
8vBYLHhkYyPn1knE4ortQExWbBHOjb4Py7zpavuQj9zhbOZG7c+Ef4T2PWcYzJiM8hxr1n/hhOVh
UjxLY5ktqLzUllbxL2vIb/bGTM8pH+c4Pwf3AsWtnb31lQliZyUsbAqIPEdIXqOREo4zlbwa0gI7
M1Diqvg+CF4Ur7BpKhLjF2EEwGbYVg3tTQHE1yUpQAkGGuu/9PUQz+8Q9FqZfy1EdZIZzD6A8qnq
j8yOPGaQN9ahjE+Uz75PSeJLJLsl+3IKYt8HvqmxsOFtcjK9796TfICyZq5w+6QIPwfq1cL2iQ4g
89JSP5qIGY6jEb/tuVUS5uyiAUto4BXaTJMNl/hKFCHUx0viTDiPVfe+BVdP83l6XnFYQdqPHrTu
9AJo3ddxlt5oawuD6eg1x/N77hsmHgMAVnvBcTgrIJVOKILslzTmcGx1CZOOXWOqIn+9ispylC6J
qU4mO/ZVQTuEeBX5Kkfv+EkTQNT9WUmNtgF62h2zy/P16CIoE+dwwrN/kPjGcZq1ig+0YXkGCcnF
17mFZ/Ey7UVTKmmeKp0D9XgUi8Mdz+1C7xoySs0KnAhwIRX23XMCFjBdvSoSqGq7OMv2bHxnHPiE
wLRQ1KSdK5xc6fMCdMOTguHbDIpVAVUvd7PEU4rK82YXY6ywdN7G4Xylom63mEPEgkbfppwav9hp
II0O++siA0Hb2CxgYNOzsXeFyIxZmJmBwvPk4UwRcq6yUQjpbQ9jGgGrjyytdOlnIpCUtWFL4dxw
KvPiLk+aJc2yrGMYHgLGYVG9XUQ3DfTtNAcM2lUTU6DDfXtmBGjbCccINf2g3muSEn9pvqX3jIJJ
Hp9z4CY4JE+4ctAGl8QKzW/QkNbqRQrL77KyZS4qGzub9XIGn12KE0btnRNquJWJFeOulSD3DLmr
RB93yaZtz1uTwwsrWP+FtXZ0lRAWt7cfAWMwZ/fyOAbypPRGZnwkxsvcvN9YWRJAwCs45/QHfn7Y
I6uBGFS8hjGs0BPPN6mYNZ9nOqoDqBw5F8QfDwpgcr/YHX8Lr3fkos6TGT4/VvHamngRQeW+MWe4
bSq9esWLHVA9/motfFpjmgYpwf+BeEPeqvx92YPvKxI/qxKORkACdOHI+7ic4YVsGlzFXf4SXSBu
cw0w4vkiwSapSFtB3Y+bbMotHt1nluPgbnCfDhUr3hfCs+jIDi2Api6MTHgO0ysaZhXGUUsw3xLT
Ric3GMfXwo+JUejRkx8UblBsq1CP7aCeNk43B3M5VI5OjrSdqv+TBV4S9tXDuRtR2hNwz/oYxhEe
5gjmMJaS82c+h+1BQ8ytRbL/nom98TnUjwX/VnF52XiUwfm5fajL0YHxXHMK9nlqrXhA+OQbmydH
gQP6ekIj3eJSbuaHOntC/z64zK/BiS/0ycEzjtxuD4vOHaCrIlTdet2WGp8mCdOrSy8wkdOkCInD
TJw4mLibWvwRsx1ffthMUcW3ebOeiSEYPZ59ik1ZWsqEHLZF4te0dRLTjQAKh1YT4nQhjQoGN4oa
NSicFSeXzqYpp6EM/cnXlrK6gQ1LpDMSSAhYkwIVLH/XVP5XTodc2cN2beBsyIp3idx5TKiFqHrs
0Z2mmk8C0uxjiJpOU+LTeaU3YRYpB6VJWg4z9AV05PNBTtptCEHCUhONJYVgIxQSDUTf/gd37sRz
8X8kDF7rQgNeOtEgUfaxZE31WZHSukl7YOLar8rkI9xr5koQMEmlOjChwt9dUw/UNEn8XV0tqDju
2pAZ37osUMceRTQmqgrvxbOAIwAAoYYzbamD3qPT4y9WEKeSTHRKtLgL9fQOqayMMaliyzHMVc0v
RI+wd9ShuqDaurOO+gnn8PZxw114V9NFbyZEsOlaRezYQJ5EUKOAflKPyva6+Z12Acm+B5XH5O4w
2QIfJ5QdKcObJHS52QKTXMgjLZdjK47P28fqdagJYE7qVuOApl8o7AYs+rmaFO1Dy8XmDgH8UPRl
oWTB3+lgFS6+H3GR+dMWMppU1Zx/SFVVHPamr6Hh8r4M7j/shM4XVcrt80ruxdt4IS1lvYHwKNsE
xQT3iwMVty8BEjchyiNDMJKXXnohUNLGI3eV9NKEbNjYVF1uocGt0oMIpzcn2/+usLuTWUPDtGuX
N6o2dNUZcOyGwSeiX9kG1TeFvG1jlhQ9gJHvile4vT5QbIM9U+5s6i/HzjWUvunYwBdzxqs9a4zM
sAzCMbDDE27Ck4szr+pvFH7BxGFgXbmWAcUbW0zEVeEVaYxgDHtC8ToZUUf0yXJEeRYO2YphxBls
bbFAlayDDdDpvgLxS5pXVTLSCYW9Ft7DL4ecIDR9YQ+xpRRMfGVoPeGRZJQuQRrayXo+WHC1L5ic
MWy/UK44TH6l6+LAGCBbGYlUzNbc4i1jAiv5qStmmP+jnlW6YY4QGagM2/eG5ju3IbcvKnaFJMKO
v0QaaxxipLEkOndxHDk6pX5ob/KsUpSwcRYUcl3brI0VkxUSKPtF4lWYDxKDegX5PRmbuCvHAYlI
/oYmo/KyiknGxsBPbiZ1fzOVMxM9Al8eTxITYuGlzGXHZN7NDXHazHPpQlwKpDz7f2Yd9l3XA/cD
Hn8gWTvVQSgM526zHB8+T6S64doM7d764c7KcpJ8v+jq6VfMoQOpk3D5scMFIM7+ZC5r61er8nnI
nKNK0dabEKGh/xWENXwkGnrLW4B8jT7ATvuX0o7W9h9U84W6W1O3mkubVXRYR0eEaS1B2s6pXXaf
PEiw+//L+lw1irmr9jZ7GhITXmvsj6ixYwVxF47bCVA4oZv5WTp2c9hMWEiGCZQlRyGeomacq++4
ZC+WG5QD2v2MPvRzFoYP9n/XutM6hpsle/e7wFw0lMtdPnjMqvXza4KI+ohauFI8uvtYtmuzoC9V
4/9+FA0BlKhDYZCa02dfAWWy0I6hylc3+0M3hFYoq8yoV/6rSdSAJSwUcvvzdl/CCee3Y/ydQYBs
9AnlifBlmdC0ixQmU/edYTX9ZxxKhFiBtQQaqHCrwT7yvNStcAWElxEJtohy6SR26Qmv+LY4b7LE
W/C3K9B1rVU/mcdSHQ8f5TDMqNgSLRNFDaG1exdw0OQtUD7DnfM0w6Mr3JlX9rWf42ZYuokH3AIq
e1xKq4oGhA3VULpbAp0QHav+celtt2H2Tv2kI3dV/q7xH+A0GZ1/kG9WoLADcdIO/48Lkx2MMzAi
987QEbMviTeGAe+hTBeS5tduq9sfWsgeN4ejbY0NTHXFugdJNdt/gsjo85htuiodmYzYSQUF6UbF
cmCUcgfdSKyrLr9uJqYZ1lvK3xRISdi/hiQUkFQXQkImJ22Kcygt+de07NfrT0t9uHvZnwhEzveH
YHu5D13JGAbM42ZoWP2VwC3sHsBgMaXpPymkm+t/wWzrYLxESWiPlk2SPNl/+mZph3iy3fZogVlk
TelUJUmq+m3mJqa5AsOvCwv/4ENd5LjXoZsQTLfLlXkHS1fMoImMKV1HOteoNLNttSrpZNAtLy04
ro67/ZByZJuaQebdZSYJ47b1qhXeRJ5sNXn0BePYmmMNAKp8HlpVNbqhlg7RQNGuLYYlvlm+E11f
yTQjPq8bNaEtAmPncJSnT6AKE2xrxTFrHpghnFsk+wT297jfprTJbz6KWZdqTPlgiQ3REbbYYInW
3nOE15TlK+OX4eSFDmNKE3J3+v1bbOUc8Z1gre5nNs7oG4EDTMx7F5TVZFDvaAZtY/s6aszyFKkv
v1PhuUqUmIfRTv0ozQeI3dfcdIzDdu/ujXEQw3X1+dMvWVPfwQ1dGq/hVSWMVlv6HC/YX5YgMWuR
UaQQ/U5Xa5h+qb8oiZlmToGpv4QS8gHnWfYbWZdjCUD1naJ3vDrVttbpz8rBzLn7MCfsHb66Q6oY
05BLF0MBT5duUNGYyqp97wSYreoA0wxMOgaO2U+pkyMN35wqZ1TXqGnx5PpOTeeB2OxtKGDf/NVk
Oak8a0nHM5qSL+i8vWMknNnNhkju0w2g3tXiT/t3Of64ujiwBxy4j4CTiXHTXMg5rYWxFLelYbnb
ZUxsDTvFFRNL8dvjKhBuaTTfPlbKFPqF44SEKYxLR8csqxsc1zIAG+51ZoxJeVGwSGx0T1oz0HDy
eg7ajqujrP7du6QGAyCpvBW/l4kBHc2VCo2/mSvhBCPB4JXH2astvrDEb3F/35BlPZaiqshS/pXJ
/R6XapiP+q6gfjCarjyneu9QztQ1SOLREylY7i78H+s9kHJACxaqHx0eGpIGaGkdmuYD84Qn6FBQ
LWEOTG7DBNYzEa0xZ9QLTD2t6y35O5mNLKBpYsxtkF/VHOeXetD9mmlu+MIYIRwCnyZ0FhW81KAt
R99eHVecTTYPCK5KD7NDQBopPrOo6j/Ngw5Mx4g2oyK91enKToU6Y/5HIfdTEM+qmNCjQ0iomKkC
Elj8u9doURXKHmcmxMvAWTfUfdeHE3AO8f+zVzr1eqdo7dT+LTopw9f2eRcw0mNh+RjryNgE6Xuk
b04+B/ljIvqGEAchGIkbGBN8NGOyiZBj0Y2IvWqaTjh1M5Hrp/KyQRenUM75wYe/zgrz+T72OkzF
tqjmXU4rcZs7ApgHLOdw4Lu56AgJ7xx5d4ebd92+AFO2f/3fmRjpf9+4QRCCbahSNgyUr71bwWko
9qXs9Bp9RGelNCHt02sVT9ouykXenjmt0PJ9iZ1h11+UhllFGg1zGXGUwInYB9oWKW+k/xO3acmv
GSCH/c4Yac6wJqEXC6aiM7oC3Rij3zxcr5lARcKMTNGWxoQT7FvN34DMAkg1DQfkuKPn782DMlT4
Uu2vkpv3rD2HOY1G2LBFGe2/begi4GeyKtV3SirqnozGQeLBTWCth0HRxvFpCyXYUPyOaa1tYYYK
SeoaSvlHpd8oP9JNnelZu/vvWr4V04T7VKpJlhZonAGVe2p+SWJmcwFG8RKAgu7b5iu+kV0MsPgI
4MgBWDjpM3zL3d5HcnuSV1ERdYG1nvbdZiPzQCKT7ShsEPc4TFeVH/PL9sGO5I589KVNC5y9xx1I
OKdq9h8zhwzRcfvqsmLHC3EalYAwLxWNighVpvM/lSHgTB5gy4ONIQwRQfBUhX1OXcP9x3t+A55Y
yXeSYEYUkHY23j45Ddz34jTCREP8XNEzInM2n+xWoR8JlkDbWhyim244AfhERJnl5mupEFK5LILV
i+HJHJZnm/7bgDsuMESWj0eXjMaUWi9TGFGI55u57k62321z/cBaPfjUmKFini1mZV2Uy/5Qx7di
GVO2xB1yonKE8CuqVRxzPLbx6bf5gGRIOstmCA+4nAAFso7pz1SFUjIp/gdBVvt7xiuMYFMstGca
t9FTUiBVG652BbPIyCTbDBjxLV7iPW59uVl1tE5eHpM97jgSVbhqshBiBcmtHx+UHuaYIfZ9RbCH
ocDfNPlg3NyTpBVFBpMMy0wvn1Pa4okUIgBzvTNOzzClkGxjFMQKKOzshfOl07UjqmOzfN/kZMra
/T80BSbWp8eMDRiwFMZV53AT01d1HI+VejRjjl46trY85Tc1fTI9FFgZ32VkNblLixn1nIqr/BBR
BG5yR0uHwXuT7c/RgvXnqeFFt3REtwuwEQyhFgsTOCHjJpO9foqsGG9g1HGfhQAEpSkh4dfgzNJz
lYga1im9PiFHz5txcZCHRpcDFhpInmnFfZBTcJSueFRgeoXF2l3fPP1DPm1ZvlW5ZjcH7rHJ6NgH
7WIiD3UoyykU/A+l/qWwtGjhu9/WP6IWt880cx/4/M67AuqAjjlbItoHg1r7WLpGd+5bFdf3qvU4
OGMkRJx6jPcElxO5/t579NAfrFLvNVbFC6FNQmH/MYkK8fBbTkHpxVE52I5eXsH+S1/OR4c9x0g3
SEaRGBSD8+n8y13kStZPfF2WtVlblX4T/c67C3vz2SgqlFMiknxPI774SlGHRn7Sa8w1YGLaFgS6
0pjvoUAX44ixW3AtOpAWfBbdU2BUvgcGOl6pOdT71EBLstYvYjlWBkPWat0z5jO1uER9K+ZRCLzs
lxICqj3AnllQRd0rXVIpHWBh6WZaDDiwsN5ZpmVfdpm1j/unlfWjgfVaLkahqJY5TNzqofEhYnJ8
DlLF14SAGasSlh3JYrBWNeVZqqT67meSHKy+GbgLR3jX1fNTn2gFQOHIeIxTESzRdeXWQhfQMGAU
H5VwWa1D8DmWxKd+LXel4xVDS5VZqqf+1yL0NoOh8XVBIQwh21p4yyFoOyT4ZkqesnU4X5cW1FQE
qXOHhAIWycLpnsBE55ipzYoBYZSc/jWxtIM7qztuLBYDaaRRj8rxnLNWLrvdO4CtmkEBpFyPrQKo
RemwEMRRuuW0UsMnF8SREAQ1H6G64BccBjzaDN28MmVCN2dRC+1cDELjaru4a0AmfYPfIagqko3R
zP2QOQDa2R5MTtBkipIIcj3WKDeDwJ69Hte6Rag/KWR21zRAjpe1L5gXqQpZEbayrTW1v9SM+oYT
+c5DBiuWhNHLFOuj8sSIb9fB6bLTpSxcd2mBK41y3q1XFmxmcNQ9NwrXeV/4EXij7aTlLPni602E
XOxlkziDtHadj9ng3yRYhB+0iFUQf6BPFFDz7vJM5d4BPFc4I9oBMD45q/9uF8V0nChOrXnjejRf
GFKIOMbev5aHyfjKXmS7TCfVrt+qDTq33Uf2PeCRtyPQVdjcmDtPbOUsZMjKgn4Xlm2SuafnbdQl
hYQIQBXMWy10QNge4m9pwEwckFcT+/aDkrw4tZWnCR6g5fyNm0smrGDEY59ShKgt8pEAPEYEC7vs
5swbRaX84zF+gItFU4tPINNXNyFL5zCeiaDcDrGSo9BlMwAmlW6v5jgc68sl3um9jBLEc77JLnQj
kV84b4v7IaBDL+Q1/oJLJ+FavLFiZ0ymO523Jz0SPoKn1BfxUPGma4HDpW36To4cyvxeHhKCltsa
m9WKjELY5YplxAAzikd1WcneP8OR11d99oeAZNa51EjoYrj+lVIjuQOWpiy7Lx16fk795Y3iQl2j
zOLdBENWrfYDIGFzvcNzMMVMWM3qhvFRjjfCfASgCWYnNQ6q0N3CPwREkY6v+XPzF3XV4rdVPQXk
DTVkWTGcbwJ0JP7fbOQxoSo+aV7/tZuG6KolqGl6WGbxFdT9tX8Rvi5RazQ2LTLwJbgfq6qVwEqQ
c33AtCK1V2lSVwQTDjQGbJzQp2mDC6mYcSrYCd0dwDoN2i9cuD4vwH6zc8SEteDzujHvyT9yJb3H
P0hmkhuKYFf+ovSdkuyclSmOfcr8MGuvAm0QBvSKzvKMLUTjKmpzEguxFXca6aB7ZCx0bMBHFAnp
3la458alHgCQllQ/b3c0BvI8hZ9mvWXqnisK0XXDxs+m6B+bKGK/70dze4qFcvLk5B8lNOWU1grG
uGt5+DUJvo32LenWvcQrmBcAn99OeGfJM4IyJohccd5V/Fx2B7Enb+0eZAR8iqsWwrvUIg3UGJhC
Yz5drGcUqXuMoHqOpMtubf9ip4qcR4vVwq4QbvVJ7P0HO3j+q0YPn8pzJtg7OkkrS7S15gUqzyPl
Mu+FNguMr4uh4aWXsPJttnuYkXMOFa0e8sWN/6DWLP6BATlf3VoKBj8eoeN3HT8Tji2gijMwZXf2
P3kURcItlL84nbNGmW8LCB/U0akaSLkgHBpCTkvGBYFQsNdR/SdKtvYKQyLbSNPI0OLcn0MGjSGj
sVN+2KApzLkdvbkBLg0RCc1lB0H4Ltsx9x65Sv7LLH05dLQjH2F47xFPBHN3yP3GJOk6HCKPbhXO
0ae3zfiRqxDND0r3BcA4UaKMKq0JOsWyU+CSgiRpv37XpblXOlqNfLzuz8eQMavbRDNkrLFqqilG
x23IZ5r4u3f4VfFQRcYW866N3j5/2AFnPdgEPcpVSkX+uaupSSmIwY9I5jOko7LSQpQHdTkW3DzU
0Z0lP8kd4gr4FRBOhZbsjUb3SvHFxq5sg7EHRAIn5osdbtA6i3ndXQ9DRFthq55NcC4gaHVjuXD9
Av06RsZS4t/oMkeG1TK5d78jMDcYFNtvk7Xw85S/t7/lHQoxf2aROgwe8+paW5MleQKSWDXxGLnE
Y+iWj79IKB9NdYbzOZzSIbSLlTKq/HVYAXSQVpRTEAyU5pUtbXYv2yscDRzNNZPQzVU7Wz8P2UEU
Njfay8gOB0dkea9wu7+zHyULddpQua9c3np8VaN4qMDm9EVVe//dmzS1TizEni3Y6yhl++KDX8BP
GvpGVeAKPfgmrce/mao7oUdJfHCpYyUlzQpBNGQHb47Z3m/PiQJrON0+9wJddEr8oyDvN1JPGuAv
kyvtF6IJShVcp3HhXjct6C58212kDQRGJNDWSw1fxBCuD7N+ynaNLPLpGf9M99XLtDz1f8WiakAJ
l2rR36Ur4hb2ByBMPi5WM/NcgUv5r5/XmQad1lK6+IJY9S3/563vLNHXJqBCl9EK95XvMKuwzxCQ
3RSkaOPv5fEPdxv5suJlkZV5Qf+79D1z8L7gFu40DmGeZepNLiFeIZl8Rwf2EwtQb9NbrlFbLNqZ
/qrVLa0jvVDTcSXNcA2mo/Lugx0Jwjg8Gv3fcZp9811cw3vIi0r9LnlkWa7e9MHoh4u1AS4qrIv3
0+A+OuNKUyII6miQVSNVtkGqwN3pSSoSytH0gMSzqe3RIiEQDqJlLl+fZEGPob9UsS1kbI2Tg9mL
0XnMjT90zIG9CUFdisw135vlaRcGGd5STOyjhwTVfjM4etNsp141pL38UDqiTepOJoO0r+2FkUIV
9jf2e9V1/1j4r27G9lQgyuYka3GCOXEvRWrMn1jlY7wfgyPO0cNAgY6LSh/pDZM9dfQiXMDRoDzY
WuzRYooZUmNijwS0umD3l+SJYA2n7im4qqS8u8CvAVD1ehBZzvHjMAFdMDifGivJYkAkNmCZI6/S
ZyW1hDFC4Ty5l+54Tg7fJgIBcRhynrloEUTGaOZqof9oj7TRJ3SZ80rxjKRTgW8hVuYfUQARbGXz
X5oc340AmautlrxO6YWEwn6ktZjHy/8w7yniZQRZNKSDB6/SvVDj+OJYsjFp9XL/7NA/E2QnkQm8
Hxhh6hkQKmdtGBpXC++LCuOA+856HI7vcVLH7QZDiA3qoBKMCw5IcqhuPwmlsr7WO94SFGwzixBw
JJPAzaeKEUfKFUWvNpZU/o90CraRktuJ/ZIsNtwGkqa0hoRgvkSqa1Llo1oS6gd9vQxqpvfvAHL4
ULzeCyDMirkSmDuPuvoYdZTAQfHkr7yLjWBgPWN3vLgQLoc/kulR7szfEzS0cyyKH2wVojAOHp2c
cl4us64+Dp8S+VRaI+jAXlspu/ORGwWeDdcID4Ur3+jEFZqX5vrFDmO7YMeARzHjJxQrhXK+6zrU
a150nd2QVSN9rp8GuWebC2yszAF6ql7OktiE/gKaIVSJWnPlIid01Qn6T7artgXyD7tOHpmZMtTo
EuiRCjBKho8FsuzrlvRiOIv8bvrLhhfXtdBASRWA9AiPPn5RbEV7KYgmh7Kpldfk6T0WXJCoTVrv
tWoQouMQMEFB88Mogng/MxcM92lCTpd0f/u85eWJSdI2z8Oo9pt4elm69E7qBc8sXJ9hqR53XjV5
eYxNSg/wuwZI/rulbFqo2Lm4yVG6NwfTqMzzhccD2WS7RHc7X5Jfkz0ss2IEmXSFnC7GV3x9UYNl
4mkTN52NlD4Bjwh+Oc3/wIONBcXDKu76cI7NQaYTd0KzHFHLmLj8eELzTSEt4hW4Nbv7vksg/Dn3
viym2Yy1PXT41UpKEseu0RrbqhJU54S4NFJPMlfMuu27zO5NzjgNcadU/hoPhjAtePCe6gUk8tCo
0bMsxAuE8DKzo7QdGtapYS6p6JkKCiVReoRgB5xzmbb6SswHXsu8l2ht0n47l68SLVk8bn7MPW4J
kqxbw5XmKHl/CcYCqnMpoinrWVaB1ZAnU9BQoZusK9w0DaSIgok0qfeVaAQi2fY9fyJu2FIV0TG2
L7VWtsyWXPWbBBuzNpG7h42gKjXwmqTd4I9oWhB66G+3aF6mu5CTwO3pDxC40DpqArG6CQZknzNH
otVlI1vd9LS66vvFglWvjc5zF6H08JisoRJkvaHUX3xEY4Dx4oyWAz3N7VI/Jiv86uAIjkhNUgEt
4MzoiF1gE/eCheWWo1JhoejnNqNfGFjfRX+mIGP/pbofo4E2UVPlkTBDOdGWd+Zzi3P6nMqgIVHp
Vxbt0F8CEDdPW4rMTDA6X0t5KYA3V+fSswJ92wqCVyIs6zyy00w0z2kKjXpFjgVJP3/Ze3DlAL7M
HIFe2YyVf7iSZbM1booSp7Oifw6CFLnTtrT21ABGnT19kaJHhS7bRA/Xicvjf/U8ebJnFqWO/KwG
yLmTZ3n+ecEGl+Pnr8O43ecSyJ04EcAOC8T0FMNOGHQA2ukaqrTK5VcpJet1/P4H8KCFEEH3BgYx
e2NlDxavA3p2/b/iKZOmjhOfbUav4pHwiHjzrKue3e1X74EgYQCUbRfsUYffdH6aJtJ4G6QgWD6T
NZDXhUypQwddnbLjyxJUOpwawN11/p2OIpYhSV6rxpKBo8M0+2F63zsdmRfWSVzJ4XVXKV1d1fXL
t3sJ1HqdkeZF0jsSVC/ffzovN2XUudNVWUfuvHsv36btBkAxspTEzietHGpE9cKnzXmfcQAbKnH9
UDnHWZg3VjumenbTpOvYL9h8fO9pD/s5gti+rFoMZkWXEj20XJ4+m1DM3SzUq5CbHry+lvfae/gI
+1ORkQMfHgNOj0cMV4W6uVNrogEVZlVUzEEOk3LFHaRHXJaKuz4HPAhUTjw3pun1ioSVS7yoPgBL
VqMXOoTa69lf+vNToNPbSBPNlNF80TdoRKXq+fyV9qvb8jaDu0Y5ntpGcvNeAo7AUXln9gbBOQEz
74IUsWGeZTtYmJZnaFGy4k9/AXpg0xz56dHm8B0Inqhq9SIVwfa6OkMELt1k9AYx0587gmLoqxZb
6GMOvZTspNz5vJtGB4vgbg95crOpLU1WmKv+1i2Z5Gnjkip7BHaZCW6HSMLi3PebF3gIqnkE8Rna
o9T2fNrVbo0Q0ND6vIPBlc2BgYEhjIALggSsj+jaZh/We90e3wNyCd8e5H1jA+umSB9IPRR/AxUw
x34taZnpTJg2w8R0I8XTLwL4ei0wLFNLlfBIuY2au1LCQfO7vZxmHbjkMGy3Yo1OD7u18jFJb+QL
drhIo2WktVIR6bf2qO0qTUZaZ3coFgLNeTO2LBXsgTxbygeHGbvdKgi/BjPZUcDmHXSHcy8BSgz3
C06bgYmIm6/902U3DyFGfHZYmeXSt0EGLUutLtjf2kRAkabcY2GcHRFMSx/r5wTXWEuRY1tAoRnF
4XFQYM1xfeh1H2XYVWYu4H3amVG74lw7aqjzOLmV00fLjf715g6c8A7eeZG/XWm0X07zD89yZjzF
S2bP+/OsB+LasK17TKod7KIaczDtvkfv7c4LStZikGAr6VDoVKVPKCD8sZXbk3CrxWN8ymV64nIF
NWTaLDyIqcZiD4+Hyi6w3ZpEyjaAuIW/6FI+fuUytCerZLkcrW1/6yq1fIDfYZefwDCfkue/gcBj
MoXtE1U/Do4IZpYZGHyt6LjhhbrZX7hZetNNPU4zWJzWUQ57Bc7JF6zf5pxvfm1pEwbPE7SaAjSx
FzsoLwaPk+2gPoouo7o3Xo8LJbRgAYoOR05l7c3XT3VvS2o6wcyUVEvEsXs+hTZS+RSpZj3jKLCT
oWCfJ54j+LeXUWVPhbG5Xu1B0kbST6z8vfYKZOwZHgBwGA82Jt61B8qm2sRXEONm73bL2ijjNsK/
aVHoqfST/bEysVwXd4b8GvWMdIp8/LIITjtwCRwuu6Mv12z9TZUoatxc+DuMunHG4wcqxVqA1oN1
E2IJBop3OaPOp8cmdJrfteeDQbfVoCdG4+lCp/QOEkBP8sWtqlWFSTtmKr5AYp3cLBdj4+5g4D+p
W6h5rSnQmmISS3i8F3s9EZqaJkxArzfM3mUJiR37UT07n8/7W4WctGRrwN1tCNiQPAQQAtwuJLT7
JIxZDyLoMs2ZYqRE1AhVzNMgbeXKyG9StZ53macIKnNAmXjKc7BcunKEy6abQ3xe5Voa/VLFKvnn
08Q3uuV358PE5MrXf0bkzsWd/Gg6XGrfPjnZPZiwWx0Z/lGS2F+i8CV/q123+IGy2HoY4e23WBfA
WH8KNehOK/b87H8dnV1WUg8GjfNWz5cR228cSrkK3Kpp6unxs/xMRaboWBh9MQnj8VY1+uLW+h6i
AYrIb/7K0w+tCZrO8eJPEt2Z0e0S8AbxxtgKA21gFy8lHVMSDbesw5L39uo/l0b++jCB4JLLAy54
C67/bH4hCdrUfNuDJfoki8ju4dcG0fh73P9MkX1XIVcY0SjaRNiCCV0atKwIa4QnWLvq55cmDvtV
qc9s6nFXnHb7KNoUbBBIeXY2rXuM4tEfhxvOwDdhY30JKvZRWAg41lg9V5mWAKNQ0lAJbi+hwgth
IDsimM7X00I1AJswmyaegfKYQ3GYFPFeO/derK6WJnn8uAZv95xgbVl0owOVxPqeYC1vigu80oPp
341pOT/c5Vp0NADsimyWSuUsgNc8uYSQtXo3/xuucgnKiMYkRaSiCp2Hn3XGuPwqdZghQ3kABi8z
O7zyuHpBEtM+76wo4eI0I3oPKxiNgi7f3Y8EL8e5xJG23HXtLGjj+er4pkB3F/I785I5bqaugM0i
E1dE4dSIJyqayJAWR+nP4fCDFlyXjagfrIQ5fQsL4HpPjK7axcAHKZVU7OPSI0pyPizRsOG9TluA
SQcVkQlwCxEXvbqzDSEX6xUYbw33YC/CqvEm8xmlFHOUo/LSaieILIfXtx1VFVk1P00MzyBNqkY2
FJLT1vrYQwCU1hMnrMKu/VdKVFqITCVwkDCvB/m+bx7mieFLItOvwBHW12PCFFECAroX/1vAZVt0
Szo31ObBuRk2bVxc/qL5JADUdue3dU5XwG3jRnGNQKaZpPW9T6kaI3ktplMbh/1jZ1vqqNAp3SMp
TIif4RR3Lvj6XXk7pvcjtd/qaBi9V08tOsjER1xgkYUZ0FEcWpxu9nm541JkSsMB8d2d5n2kc+Hq
+Vxqqnw+W8v8rTRabXfUgTtHVVzeHD0BZXW1WyRQ9OYF3z8ZCcJAAwm5TLmjJH4i8iEugGGgYTYg
Hs8nIL7NoiVR2N0nvmMWkmDkwSAcLXQNfWCU29qxP0xa9QVVlEKeR/FlIxzrAfI/fcAJIM4DYE9A
weFjTtbUM6mtC0ytxUZGKcp+xj1YrzsG9KuHha7mBp7Ok+UyS999q2Gt1M5IyYidcuk8hCZHOpqT
rmrdfdVcg51uIun3yBY5hFcWyYEwV2d0PY8a6JJ3/F/ZQQC9jeUA1L9KkUH8V4w4UYmBE8Slvpz3
qbvAR6eA2cHnP82gr+uQPoOFlqzJjVMJ4sroLnDYE80IIQvqR/g8shNVqu4XXMT3dMlSdjIgW9rC
Cjg4mTZjON5h5Nxn8yYokjI3F9LgE/bDWiQkja0NfXTioRj3sUaBRVOYcVn504QJGGY/ZwWhS0i0
MPbyYA2ATIzmpNTWylZGUN1KANhilBiL5npiE/igxP8Hz5lXw9Hfze+F0nyuwNrDeywllf52RrzO
IT4ZqbbmiIRKZaVJBc8QltEM5o6z9MiS1OEgzDzG67pOTZkpq8vGsIRB5RVLhym/M2ueAAkyP/w7
T13A8zreYlznzwW2ZoqN6xo/ePzNlK+mSmnIicoNkdor2E+67CRRFXnp0egPzzO+L769ty5c3WJ1
jqm7SUoDWTlQ3uRRlDKvNMQbWQ7N0+tVfWbdd9XhYT7RneMaFXOPDx/TDN9QvCy2fezuRulybLq5
CLL8SAoa7dABNStS4Vgrl4wUukAbHMleNfgjJsuDbgVPcPzIbqQfPHlTTESdV9z8Jn55R6IwfXtq
onTLNpzzVw5pUdEV6S9XSt4TlrMAHglFwxqYyLyXNhgGz3KIpm9Y2lXdIDCQQmzHMx4BuedCFlJf
ol0n3umBE/Sd4kilDEozYqwJURdn8lLaImZzOIdudfieP3EzfUYjobeX1ldRQzQl8B2Q1SGKD6wy
3A2Gq00BkxMLyp2++y7areKIzlL2PfXc0dnfN0puU/nQ2S4Fxn0ClI1dcLMC4XJbFs3AeqyIWa3o
ZZm4s/TzNacYHOaZLRoNsEbXjUKWD0XMpfyotYDhi1+VxCxB/2xEpzwAGGpFPrsXW3Wd3A8k9hJN
rjHDewk1/MZIB8CN99Gl55OVr3mgYM9a3+9AGDeLTLGaQqUzn0TJ+QrlTqVzaW0cCuFokfLalozF
jZM9wDixuHBhDyYlAzDUXHt9CXifUcTN8nljMXj/ix4FkuabgSUgDeIIEKma9r+tT8hmSQVzaFgO
sixF7eBwIS+LjdQHqjqH65injqeFwU1pJxUzR1sqsD4P62BVIjI1IeUs90uYf8Z+apTcz3FG6qoR
0L/yltEtiNBDD7r76jkhOuP4IwNmK1duEfEsL0cBYfwph+CN3sv10wtsMdqHXvtWCSi5J3hqcNaN
VDZKqM4BMGeismDfqmD/e7dICNrDG+rmUE0JFI5B+HLBSbDTJu1nYJXkDepA4RADJMRoKT1Bf/mY
IefbeX36b7Airg0vxLKWf4Hwed6rfM6d2aV0N7OaK1CZiSaYDE3wDflp2FwopS7RhPUvEVerl9Jb
buS/SAmcOWfO0503NieHpbHiuKbFqztujiw4Dne5SNe59igw5UrhVd8jYjJzWpLfHMPvO21fxex6
x5u4t36AMAbApHB4Ks3wm9rSzvZgm0CfRfLulcRRH7Evr9Nm7ELYp4FF3qL19j9kUmjPQ2cpPjoG
xvP6bPahwl2MdwEIWV5vIcEDi1NiUj14747TqCbHkFUchvVrBItbygTjdPS/a1CQ76zpbiWfi2LI
2f+kE6wBdRVGo1hzQC9a1nmC/+823FZLhOcxBkL+GYWeX4hFr7kba+59hZH36qgMHx3xGsQC/ezb
UfARRhTBvovdBn0VK+gz9EtdOjoecOcs0XQuOM3BYVF+J9SolbCCK6PX10qc3U9/BmLPhmx+SFQi
AUX54ccCsq+szEeTovRKDTJ+l9iKRD5zHfMiwRWoPeJFbNgsRNWwa13l0XWUlpyMqsEFXrJupUmq
QhqDypE7nmEK5WBXq2P+yJUeU92i/An9CZT55P+75QWRxkfaLhPVTixGHLbRgcVjCbzV/ACWXD8d
yAGvXhBytktdTPUPWCBVlSlBJjoB/5i1VFAOkdzAjDZBiTj8Q2Bzrzwet30G4ZphCDWtHV7GOOZh
3+9y7qXvb48cv14pauFemWAkoKgqk6HWXEt5Cgl5duoJnb0hTG1YN7camYEMqqWfPI+JFukwMeA1
Iv2zAy+s4CP67UEr7eHnZFRsONiHOVzddbTy2j6PeK11Uwq6vLpsa93x9AMN86QaN3YoNhCAhpiL
6J8UVTHsL0HLTA4lpxa1W+kT2se4lJ9kOIcMC1UbguwFZ9R5z4O1PzQY19cSQtZz/3QOmOkGXB6w
IcTvLP9x0NB/8GzqeXX/LBFViAiih4PNpy70kElIWdjk3//Bl+52x52WKO1mnZE+fczThZJ4QI21
y83eXQUP0GhKF3D4uV6qLfoGTBDGYvgCx4JZ8qZQaNIXyhbSqSt6ypC6UsqQxbxuIMpfLAefMtKx
HyeRvURk4E6LwitRQnnkpQO/zpe7E0Le6di/a3+XwUjm/4wDyB8jTF3LZpEC85brsLQSjBcG62Gs
4qPF245UITjGfnPWyod08iRkoSuJhR8Ac/rok72quAyXNPt2uScJT0TfOlR+T7+VQDZuMRm2JoqQ
TeTXatPv+fY/6dMq+JUsR9a8ZbOlQQGwd7u2N6RLfo54k/02z32ui4F4CIvzDTdQGlMTdbgzh0IK
eAC9FC+wzFXwQTU7FJAQylel3KMiFg8X1oFou9taOPhluCjU/akMgM/LzyL/y3cWaeIzY6/1YUTF
H2TXA1pEajweZIBGQu7ep55npi5nBPdyCvyAfgGYPbDgUou4ToJ+Eu2/SD9Uo8MOm+Iu5Ow9K1k0
0bfN7abKadWEmtZZCQZ2X5pxURMo6cW6Paqq3YwzTgGS6U36ZI12RRKcSTnff+Ajoe4gXoWdwf0m
S8uS6q1SnbqUCSiVOI6Jn9e4pjNs/UqLohtkRaYAVSV7Wq9HM7H1FV0setzW1bJ6CfZxvmDOlYQe
yoOXLj9eynjJYQpsIrY2NJYHRP0oKBeX9JOLTIxG3mI3b4YB7rKgwclDKxtSoeaQT4czUchScaxU
BjHe5YqfC9wvzZSmYsVG401i45LIRg4VmLm0XCvE/B/qqJcq4Fj9r2aveJjvQ8QUtUMyqnf8CxYc
Xd714s0Pk+1q3tq8AaJcqebZ1UJNGsLiHKH62JL3L3AeCEd2wAK1c+Q+fEOcre2U/P3mR93BYY6E
7tQPs8KAmrT+pwwRMvzK6dOG1YEMUvUw+Fyi2kaZZBzNLaN8pBPA8q/nyUG/WK8AO3clq+JO6BiN
hLloS4Qj5IDnJyyZCPnroKyQmUOiJsVnfMMSb/dBxZZuc/5MR/e59vJeNXmytOLks5d6k6XlcYHo
ZZdq3TxK6k01I7+aXlHBbjkEA3TH/IctdYe5G0loxuvGEZsiCZA2UGlLYsyezqeM06jRpaOxjTrm
sd2go+lIZKJvVS5PyhEHNlxEWT/231KafdZjqEfZoQWAYpZ+X1Hy19EvN75uCZyexuM83Y5XdQ4e
y872ZJD9y4aUeciQwefRhAqjuZaXxD7FE3geX2k+5D/41179OzHY3iG6h5WLTEoiots9PPiKAJ2S
XLNdX/j6vMu4ArzlaKEnZIuKg63xmSgFsEyK9vvwOL0vbmy0RjDc1HiNE6Do2ZIXoOWo6xP01Xqt
3UC+Mjg8KtC5WNm+HRTlL+UX47GL/DtyhgIQRcfl4JBoU88bAVAfphOfhXVMMnkdql91myIlmt3A
jTHZtXNY52tKaisPqEliIHwWFxVHTPcMafSLvEInPK2nfiMwMzFlGDbkU+YbMbES/bh6RDAn9Unx
RaY7CppJ4EmkkH1VbrumOJV29kK434V48NDQmRJ6q6JhOLDkYJuOdNAvFGSCFMRF8GGZjQrDVXvC
dyv/B/XvyAhL+b9XpMl51MJY/j/uIG8S8Hp+YwS6l54crUH2Za2XrqTugAgFlmSPP83jzH9YdRdJ
u1/z/EYqcTycK9WNAEVbQQnSHYnSUah/8Sx2Jvi9igijlF+snvSd65jqgwhcbSaEVPL2sTD2seg2
HNrCtlijbduFfI2EWzJ1gqGlFUU+exBMcyS5tjpKw6isJ+yJsdmdBXA52skgumdgnDTlCYudFKeT
ZvvsURN58VDLUm88z4y8GlIER0z7ObDtHosgDXCIzHJhe+uZoJ89rD5L4O4wwGAAIInLAuU/Uyyq
qYX4QUM4md51Vqnk2HacJPlGbc6he0MhbTyN/+LdDTHNYUVgIJKaUEn8YtZvf5CIKsU9n+t5mcaK
1rDB5blViJL8O6Obig2u80jMd/PWUv46/5qhFsUbiJy73y2rvlzEgWsYiuGr5uH/FiGWM7P1sErM
bRkUTcq4bYAPZXRIDYF2K5Wvn2yL9BwI509qHstR3Ye6EU6ccNX6i0NrPsFE8zBLwrKkvXgdTHSK
U4b6cYxYVI7fwmKMGaj9z2RhOtn/MnoMAWiyyyFMQYtPRfN5/5TfCClB1tC5YNUHu1rSFOI5PNSl
hooP0mCHHgSXaEVcf5hg+JumQf47JtX/m+/FqJJAg5u/o+nedOMuKx0VGlPZQItp9qGU66yO/7Nl
pJ6EOSscJMSSaWIlEIclUch1yIgYccYzI1NLcuIHx0ESLHxCrhcNohWKrjoTWBjI1605+AjchOez
pZv+4MkPea9xjVRzQqqq7AfnDdE5M4Rn2uMixBPOslDtsHHr8c9TTgd+AL5gdf0dxBfxhmosK2L1
cnGXs9irp08ZHGObReDnoVoW9oqH2fttcW/6ZrLip4Kt6EF3onPHIOiT7yuT9NEl5JfojPKgSRIX
9NaCk/Nn1E2tATQ/atvxHPIGoXefkkQI3YI02BwfFpBkl/BNztueoHtEYVDwgnvSEEbp2RYaAZoL
fHyWdujNKOUv5CFROtstGgQdLLzGrr96tCmUx3CTIXkbTrV93hhQ0gYTSeM1ss/Zg9/THxH9ixkH
uDspt7yhBvNB8KO6TlKeoQh802RoU4r/P88YqRbANVaDcs3njPyA3aeUwzcdJlrNddbSEK//FSo4
vZLE7Jlvygl/PIfPkZMu72AI0wyPevdVg+hZ1+tUFQI7FAOrnTE+e1hbELbVKYSTofw7m+XNhnh9
+FyS5U4SpTeZDWI3j1R4RItshKgDJRXtEUa0IBF7LCjG74vmxq5p3UMdJ8v/D2HcoQQOEsnUDr/o
F0hHP/i0x++TinJYA+qfQHAyRGM6fcvT3BbMibfuMoHSVz3sMTVffaeTqZVn+Pq5Qlb4qGuY2BHE
7FVKg0dzxz+Inr8TTVxAtEZaeAdF3j71djNjdgXzEkJZNTJPFopQbMfVw3p3CpTo8l155FgcDw8+
mnoDPS/QRjqLw9rpSu9ZhBKub0gox1mLURlJMC41MmsxjMzTwjOudjv8jBMudKymkQW4DfV/Obbo
Sg5LiyxyBceToGOgCFg7FO7P01BPJJ1IXp3ZdiiEG8IIyM0QGdxH154GsLi0BXG/0Uqe8jgGEecX
T1mj1DdJbPlcLbiF72AIMkDqMWEhrtjt0Ck1zr/hGdy2TBCK3cDY7akowtWx5UBghjEAQqs7jfu+
8pNCb4+aUMPodWiyTWnLujjth148cLh/n+jb0iPS2U2hI3Z3dQrcuoQXjN+WdXMYa4IHQMMY/ZSF
/zPlAuB7YWhipUVkg+AejbwNn+vpa96ZnbPl4E41ShXObLbfXNjbjBXctxq5RQwRf+zDrIAmKoGS
YiI0LPfy31ANxxJ3jXEBNq/90HjoWbIp/TLLk2VyRyz4+dFfLa8I1GmDFIeRlZ6+FkoqsfCnQSrb
RqBexYdM+FwUPRvtpqzntveoy3CI65Zcwl+L3z/lupFz5Zl4EYJalw1hoGOQ/jZbD9TSSoGCiN2P
Zm9K0eVYdeezczUzQpJrNRnnTcYehtlEkJneCgdzx7vdJigX3bnwD8hsw+2NCrSgcGAbsH2BnL0i
vB0eAWoBbJp7pijXbGiBGEb+Fv0htICd50NmGevKKXzwgNcygmmPbqoqw5QS5qsAWWT0KUXXGicC
WhiiLZIK0Ug39S+ELBDLjD9phd++FOoLqovcM5YiaZcqMjMljsAAQB/UDSSYO63tWZKzNgNMMsDr
FNeVM5wfuxfMTGRoB3pBJtaSv7LG8wCmPmSL4doouDDb/MNyXiNjyC8mGIu8IJv7NSdbiIUmJZ3r
WynDYortgYW+Gh5c7zvcI6VRaeTFaE2ozvZH2O1IFrXiOppkouaVO2+iEqBIHVYQxQ3N889spBrp
Gx33tRGaQxN/C0/uXDFy9MJtnQ8yyd4090LZOlvHxHsithCA7dF5SIb5nWMIZP+V3Q/+dNZ6pRRF
TAC56l1OEPHDEuY4D+lwgZyVJHhY5xXEcS1TN0ke1vJLYo70cF9t+jb/TE1QAvEjlxOXYDvKB/w9
IAHoznxIZYKXJfqdYdWVwXxi56nih+VpecfseTZ27NwpDHhQLrpujbI3nbb4gBg+kZlcgJ9YX6vU
3FihwRFrSlGbt8O+iKeSO7/1Btkj3H5Q9LSPDWpLwoQRVHDL0y53y5VPFsInO9KENtbde8DddEtj
uQJ8GgMvI2jen244URz246wRy25LWeKYflxiTG1tN9pYzD1HjSjLccDERiheoNgfnWwg8CvtTxZg
P1rHgznE0pmsDmQlicQC4DFeK5VmhHUk+as9nr8Uvo0yIqchMbOaTYiO5Tir0L0c5jZdgz/6RSrk
kR3Lwsf1nskucIaJxi/9HnYw2Kb8kZm1el4upSbj0S4xbbCkhuCTDBsF9v8X0Xhodx343QJVZQht
BaN6o88Q+A3wsp6Y03Cd3hYqDEPht6wB397h2ejIw4slhzdhyaZG+eMajmAcbbCQf8jYndluDyDK
AdzY5dUaah9Ts3DhRdkbbpXQ5QtyHX7b12rB4j1cD/+7fVGsR8jVUmg8sy+vNUSNwXUgleHHMeUB
oEdxvEida9CDWfc00nPIf0J+kI+9sP1fB8cPF+SNTVqy8mBC09L+s4rNOflsosO+kKHKqTGMWfoN
r7ztbQRKb0zmslUUEIg6j4TWxvD2MCayJIDRQim+V+91Fkanii13LOzcJHKgcfBPLpVYyEjy50mv
eYyfe8LDisSA14e5dNXU06YWsPL2SrmcKB+l4FPwRetEnbp2ZLSsHuOOSNYw38uuUDxQi0Z7BOoK
46qlv6utRJVm6OEvDKO6mZv1fcKoISX4RIho+TUmY6Wo1O0Awhza0cPBp+U/StfxXrIvN7RS0hV+
4kDpR/lK4SnJYv5W7igs9KZ9AKpn3nxmXuYQ3/+adU0Gf3U9lpK/ueEC+7Z8+qn+/DoWV3ZuQrlS
zRY7J0Tbjz8ukupcTmm06V4VtF2RB+MSqmpXJDNxOPaKkdf4rYocaA1EvzX4bPt/DUO+DzumXyWf
N0RUoD7NJYUS5tq2SObg7Wke/LhxsIRX5scvVC8qMlkUG4h7LcwXZLxZmVnX0RU8n2IHbGkT7cPg
Wx66Xc0zl8lx/PopxgxZUAZ4yPYVU0dMKzVPKFUDRg8pIknql/GZu39Yxne9OkyHqq72djZ3jmbU
Sn6uvxyfkBj65Tn59BRlw24b5Uz4cvZseMtBf9YzUrV4OOjjOS6o185QqOYP9XIfOnCmKKWhgDzB
ncruyM+uxfBK9JLnBHvyKF1Bn/yg5ZJMAyDz8foAlXuao+Vd4TrA3ewRlpPZ2W7fvE+tR011ETCG
Sida0d1MZnQO8nfu7XY2Fr6Q04tfBqaLIO2V/cGShyQttSTmGRX+65xEX3WurplxJFhT1tzYLeLd
dXuaPyxaB1oJ6eh0Py+xSOGgbvsBP8LmoUdYHI1DW3+I9oWt595BjNukQTdKao7t/xhlHyQfnpwM
jSLj0D3+/pgRzw2S97Vc981pTXEEVk13Mzviq3in4uFx7zvstiUfIgZqlKz+9UyQRUQHVhVs6/AE
YCI8AxIphhGRrggKyt3nQlN1GDH4xaqYtjbgetIEdN9bmSlogk5vJcuPxPi500w/AtJyhZUSm7Nx
TZCfU7jz6wPTeSLsW/f3B5NWRo5XUmT4FIwX3q13cvkZhOymtTw0h+JcJHzjf9eII7iuunEQI7kk
Rn0GzBqGMdezR/sI++tFCRboEvkFUKwPi6uOU8wUpBvZCqTEDbSREnli+0ws+5UC1pV3yrAK+t3N
k56swraHtOWBpdWbyWRcviLLlFZlzNPeFvcxDMBvbnoevPelWQslycHxkmQABuYSLb5nPavkVbr5
roH+qST10XzPPdWbFCdFjNsg8i4ATcbatwlHjJ/qRNFNv3yGBM3uQm9scuJ6ojQ/lCek6D+utwWO
JKWqgzPkfBDhOWeHFNEOJyudhzplM14g+GrS5s1beLt1MUgwMUfx6+2RQK78qJLpc1/mrXNgx0tK
TL+63Jgmh4YPsxgKEQSucxqH3X+dVMVTi/80mQGlDhhxoGA3bTWUo7I7D18KoTsjGr4rlLs+8rP/
F3+UabtV/NCBBD6EaKlXLoKNQgnE+jTOgr9CSzQ5G7/ogH5KrTis4V1Qs1K5qC4/9n+H9N96qY+S
s9EhryNLWI8yN4TvTZadgbgnnZku0WFJNb1n/rZ2iQOOvrpTDmrTTttPBjvXLs5MqHaosJY41wrQ
xfHjJstqtb52cttJh9rFD4AZXC6TsXug9bEeRrwgiIt8AWNsHPSV+0xTkErlb2nzpKlLMRk2ed7I
zs3ccM9kd6K2BzclB8cIRpelni0HM8RD1amJw2MplxiEZuwnz8GgteeJMqhdv5cG+s8FMU9GUowA
vWWk8+Bsty5aFA5N5uWdsDyCNUUInlqitUbeL0QbQQ34PPz5In1lSvbOepwq/SonHxFB0Q9+geWt
j/yn53fyVOvvRFNxPpzo41LRMdrIgYZdyX1TmUwZ6kH6GQgCdnAuJq6chEaSOtqb0yfSEAfsR3mY
/qScE4655YkOmjwvJ61L/kB2yVS6igXtWzYEuo4ozwevTNJnbddtoKkWYWsTh7NIkMufAHqHYTtg
nrrUs/Ie4X9EK/efTEDeIU+qXw/TIm2U7pKXD7xUywY13mvg4WFRkDz47cEbNaxjjhJu6rIH8WHN
na7Nxq+YMEJX6N7VK/yKmhNeLL1PXw7CEoqTgAeGWDHfeGzqF8YM+IX3RFaXhiUHvEioy175FYCL
xjCX0Gato/Xk6q7l0iZY64/lLPk7Ejx+2OH1Xzhcqk9MHljkQBQOin1UDpiesPigG3m22VAigDjH
bE6VJRBGEgMhCxNQRn1u+slr4nGOxYyFnadfK4Vt46EYKkTgoez4x+81244LUz8usedZKaMXjQvt
qhPOXh7k1rzcR/QoDxNoe6JWg0NR5F+/Zka9A/lg/LS08CCOnVTfk/C4YxNVgUpwfKy5aEC1ArDK
ckSqMFcHrazpaJ49LZRfh79kT7gSIMJbSSFp5mie+Cm2ebt+hfk2fDCHJspUThxDebbBXQec1UjN
yaekGXzemVt98z+oaZJeHIqXOGy7N5TklkQaFS/kA2OVLekNln+C9gSpEIFO32Tk/gNkDnsrb42C
S//RP3L8A5ZxTD4C4dDQojyJTyAdJBQ5mNRB33kM9Y/E91K+Gi54YlyHbCmmw4mo0XQXM40Ba1Wo
SEzm/UkPiHvh9sqGMXxwMDcdOaxowCLF2odGdHw/iX87rsd+dN9aa/G24SVln2ZzayGuyJ1ElBnH
lK7+DWuFJlXwADlQMCRsOpZH7BTyIvMjIQE5Y+zYJqtdPvKbEfmvnfv5G5t0fUiUQisjZOCrjYKE
yiCfxBMsVOjmRqojVVNYhnM5RkEBTumzHiExRYSsHf9bSyrfxztcqb19ltZNTTCcAG26K8uRsHGb
0mOfucGmgHBrXdEstaL5baHEwv6R5e7HqJrjvQWgc6/rtGnektBeQzO+BkHIZAa+4t+XnuEPLi53
hQQeiU42ACUJ8SpXxt3XHXNmaFBtdIoTxV6jGg5QiAA3ffUEYf1iny6u9Cf5VNUzPR2Alx1xukeO
VH+ug+vrdzIOM/diuS0P0m1rL5P/kOwK/yK0czKnw2IlqZz99Zn3mBQNDJ0E6NJzNqGen0pN2aVM
Ih1EzzlXeyVQki7/YhDPHHmbd+nmgpu5jOIJ2cXcAJhHkxDGmF0ogMcRrq0K2wmfx1W4Mg5P1XYN
ouvejrZ9jI3nB9xLPcg5lw5giQzCVGdJo+vcq3hA/g72KLuOTO6rQk00rIRSmeuKkfLhN79+SldZ
k9e0NzIH1/5lzcyJ5ut1yqHu0EljErJA/cnHe0xPU7V+5k/IYR8Ak2qXbExp9cOe39qu+V2Mdu5r
w3RVdKuT3ClQaBHTSG7V3zJOVuvQBkceo4c1VK2qtB1EN/B/lOMwBIRy6FjK68xgXdhSnTJ0UCt9
jCLRhGsNxordWs9MT++j61/3n/2N7Uyw3XNPHmjAWezXDV5zrWBRvrAZv9CZeSW2whEaUHmJ/krh
JBMjv/FzY7pOB+B3cX57tqMjkhVuzBst9xvrPtyM4unErfPvh97hY7YxQyqYI4b7M6gVp525x5xk
BLsVLrKVgfynaHwx2Ybc9RnmYL7htWhlvbQqFWQNk8ahbbaQIg+64RYQDP7kwxm5fpLSlU3PhPoc
+VwtS44l6QshiakGDJ15va9g5xr3u7nmerwoV/dhMPYDl2JUjZck7P6eqssCuAyothXmbmqhzIRU
HLM1fNBQ/kphca46tq+37hSGFycZfwoLbo91lI7BoQDysOJdzpSDqGkW4XkQyfFmptdrWSHQVpPO
dXEkcwx+tMebyO/DVcIbBCRpid5LMxqLY4P8ez/3Za/qvGow4j2IzNHhpbgsHjIaRMA13HbW/Bsr
30ncBOr/q6JVQwKjbi8AsCQ01EaQkv4bWQBOfU20xJdeNT91mxBUyy0XzDXGEerGgR/5pg/pU99m
TyQRGTTj858dBpqe/H+toYAhkl5LjQ8IFjYjYPLm0V3cL5NkWrLM3rV7+HyNFQqlE4HHD60TbLha
HJTRPGbY0iHXeM86AH5K6mrmCQNWl2GqdGEnQ6F059+Ko3a82I/fYRd4/6AUWl1eDNurGjNxkRLM
GjOrkhu+lPRJBfE1mZP+ErOuCtqGOcXWlFnZm7HRniyo1XedAXe52zKbvF7u5oN+T2tbZe+PdnFp
3lFUeRGz81be9eGrUKeVpLGyqx43iHt/0x8mZjfYFgvYe0y0Jn+U1nGYjBEf0ro4n2SWLHyK7pl4
YLLNCWODDfaYbPd6elCzONJwowAm8J7zpCFtQ0VLpuqqBTnqpBKqKu8XbZlc5vieMzx73xJSAUOU
nJFt3Bd8yo62e4p7Ecszp2vDsNP3AorIy2z8NY8qEHfhgz1kJTqKuPqn3oGtUSBgtUUGY9IRhdrv
19bIpAOtMI1g+2W6fZBTPcMGr1eHWt94bQQp6XeCwiYhCiqSFW2yJd897i66xX0lBL3XKpUOrNww
oU0Jripm4nbEUeNZCjTncdhLBkjk4clpgA7aBc/L42NPm9SQmlVhYZf2oMIJpGVKE+ss6OOfgZBt
BnOzZ6JSHCbtdlos1W5yv6zVkKO3Q+vh8/kJejYh8lrrlNQod78svAnWKZEst4mETUdNS+vQYJUT
tfpA3SstvayMKFNpQCDh8g5Yd6usnaLnww+vAimWCde2jdFzTJ7cZt/cu6I0FEv8xiCOqMOWKM2s
JZEgZVdEpZ3nhYj8yWI089g9SL3HTwOtT80G8HRTJohE/ndDDhe/koGPy5bk8l3gvFSglqIAZRIT
T1NlU+k5V5Hw6ijPVhg0Fh96d84UU24v7lNMDdWMFAKIZukUxwOhlmEQReB4N6dUbAasP+nsfLzw
u95CO50xjdkspePzs/ZvT3OtR7lMcmCCy78kIr89yr4DwoYYLRgrGOFWVk+wWXJMmmxB89LHa+uK
ThzchhBhiTqEMtNZbmsRaH3zKs6y/MmS6hQ+yqdKNj+kHotQkyCwpXqpMjEAX8anMJRe1OikzrUg
yfgrT/KuQtL4AKCLihoe3vTpqPIpRLz8or8K/KJa10fmwHfrjq+kFcuMIf0Omcr5cofTcYgzZKcs
eeHCV2OWrrvid1SAlq/zlARv7CZqxdgrqDwRxhlPuulFXC7/TMntJzlbuFmOhUhWj2MUwuC+SIWo
4HRNRXdYV0xiNAeLiaUdNTHCoRPko9L/n2IuT1mpt2Rzc+9XzPRqk93uVu66wKrZlL/aMqXg8JCE
asDqjaz5EtxId0Bj0pbP70EPSWo9xOxgH5nWnpXXaxwO9mzlOtZLyvTwekHxHnneCLp32vjXcmfe
ahQwSraf4oP5/P2DfX2DxWDxEXEa5+8x3HVabccu34om+1xBoeNgy/AMmBBECDloA2r1Yndzyp3s
n4dRMtdpL5N04zgSwqfc/ArLZV7I/VblGsqURmj8epbYW4mQlxZ2uWjca0VHb06n95C2uFkQWDrg
OZ28zcEsLoDS7T8Agc4ERTZ7MF1iYin5QZZCob3k3n+MX2asNuLl3z0sp/34ouLuTFL9rPtYnF5d
hp4gC5f5GM8KH/qMNxzB4XHJbSwEXC96dzqrwFiKuo9cNFUCloS2JqCnXMDPoPw16u/OfMywBtRT
5FK7ZylVZQKQvmpDdLL48yqUA5Qpu6JWPHDRRXB80n37uZzSwPuqfZpBQd8n/nj50V/5TemDoWjT
J9evw9FVC1CtZXeI7iLVFU0TNBuM0T4yppKMlYImBV6VNpFC3IB1atHgvDZtAq8WaOSvthuJYxuB
rHXpL8O8cobpIpElSUO1TIzWp3qNLUC27o4SfFPjRrLp6Kepx2VMXoBiKGsUHJ+daecbxROKOVtP
c7rM6S2linYfUbgKvrBfkH+ONdsma11jxcHLN1gBVrhTIuglN11e/LtGJcacIRSYmb/hjGBJF86R
vmWYC4JaNDUXYRb0TW1XC+6g8iX5MLgri+D8m27G5IUUHDUQBcD15vfhVMPHdHtm+9h+Mv/wemrK
j3x8CJX6JnSaIssG6t2T2auv3gUt7pu2RDa/fuI2a1xSPJaDEgjY3ORJBGqJ1kHimqj6NJ9U3bMk
k2khmoJvatSjRNp8MX0WkVciE/b+D+yVB+Jn0onOHUx4Mi2Q6r+abwaOvK8TemGnS6xxUpoxz4j8
gATHH5+58bylfXrfNNFcgSefHfg7hsk382z1SZboNGscRSplXXjZtxNrQVRZMWK8NTFWjmIIy4sI
W9P7Gf49SIAXztdBqy9QTYiQQK4PPCt2bZUOLPiRcIeBLVdvPODg/vlW8JSoQ3n08PnEkuLJm8PN
PcSrta6TsuQ3GmYx5guwRmmaFObE6VXSf+Yz2OGXnMjGYrefgB+uKFayq7tcuzbQI3YngVD7+hiP
XwB/6bGVidKRILH47HsNacjKjuvAxNUs8/9LJcrN1bYwfWboTVngvfdXW1uKKqr3G+KSN15NDyu1
SuWGDPUSKA3LhTcyNUdsgxMlXMD/BJwK9pYtWm6VXcJNbolpn6X2lOrQLlBp9qokKQ9qRQe3jSX4
1b6H3H/8wfD+vcnlNNsJ9AM0BXEq+ctLl0Xysh3FPjT2QqSNRa/gpdvM7IwuNhT27/NHevdTboFR
pzyJfeyc16BTP6jtX+gmJRlgx945j2xBxLUmPLX+PbiSdRqtMUixqkGSF9zwRLZjisx0m5VJwrLC
+U0nQTNwxs9E4uOKASdyABRD9PXR67kXbLswQccrIfAF+VD5QeWI/zFhgoXIWWUg0ym6z7ABFBS3
KHMZfeNxrTVk3p5iWG2+F5c8m/K3FGnwZN1iPNfW7RFVSk4ziF0J3N9wp25sVgQMJxldKlRsRqmc
KCz5vwNZNUw3SwWiKXcwb8tPpuMPYYaHo6UhNgbY6Nc+mfozbmRmW0pdj5tCcQ4m+CgnpMbkqpD+
VZMu5QLOcn91IF17K/an5yPkyXdawNKaQ7khk8xn+v4cMVYd8lmCxY9L7sep69cDzOuyXPnARUJG
0UFF8CEQwh3CzOq9ymesevgmaUXmmruGzsfOMhb6hXBcMHrgReVktLgM7xwDZpy3wlGTLoJx/J4L
WOzRwJLPwJx/8cIQR+pQQ4X3WlVr3ecrmzcxh2tzHDqhChl5Us+9O6OUOgjvJ41dzzfMS6/9Lmsw
uEiNFnUfCJ0Fur7M7MMZXvU8TjjpmNv/jvSL0btUt7+mkV7nl4CfnpN2DhvBGMAqM2WzZWrQt1sW
jJoGCoGocOthE7vz7HGhnwfecnj71rp1evw6ZZQHMBh+0GmuiLeeaPvInJNXrMuYpE+wEJIa4UPR
/Cei3I/q5bLrXUURrS2sjBsQ/1MbpJiR9yKKMSnlxTw3bhN6zKxFBBn6xDyLJHZEG1512NDXUax8
/QCw+pCBC/Cf77WuxBEJ+BmXx/1wMVZ3FOeklAXWV02Qd9B9LEGRFnIcjIRNjd3+QOzJ9t7mhj9/
g9yxXP72aMV81PAQmgj4mo7txKK7D9nUSn0lxO7SsIm7YB6WIwASzgOrC9Wz1EexgVlPM4lG+ZKz
3qNU+l0K2xa0g4TyL6AgvhahoRmB4KWStsFWqfMc/t+x8bz5QY6giZsI25/RuXwYpBRUCvSM0VIl
ZXzqZ3C9EsWTVA01FTbptj+E2c/k2Hl1KgGVwBmFdbxvH4JoqpdPNyvHBP7no8eV5RS9ph/iQiSM
oQC2WvAvC310gBk6XUAZbR/v/YgHSbIxsbZLsqqgdVqaGEHjsSkBv003dUN+9t3vmSXjCrMAXntr
XswijQOeHjmT9lsIWC1NFHAk6FkTu7G09/Obk/4FsJaj+wz6bzXZQh8AMg4FldcTm5TtdHrEh2Gi
wvg/6HiqSSKDriFdtCZfoQ+0bS0rMzJCkDVgpViFuHwkwCAjmqtIZIc1haLPfKG52DGdiyJhwI2t
FwHdr5CNYlaHRM0YY2g7UX33Q5QvgbaiC6I8Go+RWQX/mZziTzDH6RqrOnYiWeh9jT9XLIqPe60K
ITlMSzh+id6F6EjJXSDD9bcF86LcY3xVhi6f+ffhKwSsjlCcVSrgsLpaKWQmosZY0BUsMBH6TG8t
Byjug1eV7pQfQ07AntDKv1s2qwHnqsUm20KVZwmI6tQMlWQ5psJbS5WO0F+QE8dU34LY17Eh70RJ
wKV07bD4JDHggNfVify36NQwRfC1rhjfJoVoOfB8RwlWsfwrC5vCdFrqe//zlzQiNNH5AnmDzDuV
KycnK2XVh4z45jJ1ePZ95YfVuMGkviBp5Zla4Tna2gc0oyg31wNRyzPheU2wuq3FYCITbDN6787e
bk2ZJnJCAOkh7KKje0nMsWvzuqNLgMpcA+UKaGi8wfI79Nke/CQfDkoz44hEkp9wc8ysd/tgCdz8
iy/bqeKwpRj33R/DbxXsbKRYErBK9KSBwavzCMef1x31cbYjF7ZN0YurGjcZfc4KjY6Q/xc55vEx
HgO3NdLQRuFyywxE3mvUd9NrMODhmoKkL385pOtn794HNglcqE1lHOqmJ4AyqKKQf7Pl5FpFY6Xy
C3prfr6FUvlKjpRpVeflJT5sGFyg/hJ48ll32eYBHZXrAKpxFBrjr0dLtKxzv/5w+vzi3Kt73lQI
XKzX++lVD8EDI+TKSAy3F/6i4+Ml6l7tVIqWwBnS4sopdqCQ+Jy6RDZynwTWJsBkteyyrgHUemjf
PdnZqChJvtKt2WrFcIguQRz1Vh+nkZYanJK/HZMDFNsUaL2mc0tvmdgjr6AEhK69wGCZfqhtg2Qn
lESAWxNOoIZakt6N5zK4BFHANENyZDBnb39gw5XY1kQenG9SeMPVLrPPntpT+F7fdHsSCzZvVN16
LqpxZg5wdqaGvsD6KT2hS5W+hW83f4UN5128lHmcVdjyYpGnQhbjgexZt71SpRj4VPZn8M+zy/KN
pkeiWcL0PAYiT2QrxSGf9B5XuTrAv95e1gaWVb1fkI68xIzuiY7xV0rUp9k4uyxNeKxsTebWmq4e
fk40wNGDVd5IEF6Y1dspfTe1YPiJRa3dudxFyR14BHlVj4vLKziq+U0P3/VbHftRcBG4mMQVeOhY
ZM6umZorc0c3/Y7wIg5ZcN5BmZJNoZMgV2XiyiAEEfJAGhg9hPstcB65wz73cKYMtaXuAHvtLYJ6
py5paG7Vw9caiz35o3f3i5heaejlBrXVFw1yJMr4w4YVV71VVNMR5ZXPQuud3L+OeC9eBk3VaAuF
c+wgkDGrFjieDQDV2WmsIPgJ60bzU/62TI6j/AaE+pBdY+eU7g591S6GvEyqIXP3P3+wQGTBeRwM
rVp+EODzQxmA01QXuLMV8j6fM1Vg3CTPZkomhIugQk+R1EA9MxuB7YDk2UpyzWU29pZPutDHg5SK
QSNn29zxyqhB7ytiC1aNKQFFQLzXwpmYVGeH+Rdfiw4CQa9pmfiqi3evucyxd7wQdPMsen9NHZ9b
F6Kx9nK+JwiMm+meWQvjgVRhVzaWRSGdyb/Nv0Dg2bvN0LI1gRUsjNoyPLYq5bpymHJysJGP2F3I
XKjTTnqVU8lX5JiGTpT4ZNPcBH7flyQVaJVooPF2Tmc48sUUOU33h23iZtA0WWLTFk6Q3+4OpNJJ
a1cZng4IPRMbzdRNv7AIYwDs3HcrOp+ARJ1bd8FpZ+unTYLoqdMVwhxJ7hJl05qJ32A4QO/3OBev
VR6bfcIshAZsY0u1Eskg0+EKRDY+RPaasJ+yS5qi20OFHetvZerWPxMy7Ke2TGgR8OyhbnsdS9UK
AlJd9f53Gh2piDRJHUgANk/2NHbBoweHMsBSHiUz94PUIk0sVFasyBIIPUh+yyuBPvklO1ih7WfO
esSNX7vX5Z+nF+j5Zao9tgMEyCqoG7Xt5fievAXKKlyLwMZqykU5OndGKANDQtDaP0JAx7koSjeJ
+AngN3OIX9Pvx6VTzdBzP1fW2UhlcQPR4Vp8pmpFhYZ4n/fNBXG3nLs2QRiCpS/x4tn0vDSZp+2E
QmP1QkvDa/bkaWZ+RmFpsGi8uY7XcJnCxLqwCmbzJ+CAfha9Scb0e3xY+rjcwhlkyisZKx2s1V81
Dz5SG1kcEdQH1wWVBvr0UDWOZYq1ri2uMC2zIYnbpSHttNSsE8aB296rNLCs/8bGYAgzZUHevOA4
exvOTpdfWtmaKjSru5Eh0p/eCjBRJSW/Roj0HvcncfN2IwizTJXNWoO0mnr7p8onlzobrF9pUr1O
geol9mwLoAQk9mNfoww9JQw2554YIXMV+wkVyIIr8Abn8Eq4cXjNwj96Gcvd7qoc7zskzjY8hazr
zEVbunemM6hAnlhcvk3RMvi8VZ5ukbc8uXtMh9YjMWVYVPFk3M788t9ONsBGtFAPZpczc6HxyLx3
q/lTrj6NxfTY9B9jzm1/Z6cjCL7DyhtaJ70A6uiI15CGg6o8bY8r5z3t4hyuo9pBxH/NNwjNsUc8
xSta9aSV/ReFgnQRFLbU99npXnFnrFljIos/zxS+RiA122VvIr30ethbIEDjlo5C3JxmIgC50p8R
VfbBySn0+NmpGPcg1D8wBMr8Yu38JevoUI0lshfOP0JvhQ+72x3GqjbvVHH+59VzzRIBulfFsLbA
/jbpOvjthuxFhZyB4CH/VXOHaOZVaAhBZuDHlRxX6JlCji4q0RUeKxcCG/dRb3mgp/QAOEOr2WpW
QLO05JzF9UPN7ma8rymNc/GpbpK7RxFkZrMdRC0MNS5SPDwpmiNyOBASzBmAdlyakAkBpsiLUfH4
xWA1esTGaq4wTuTKR36D/C2NxBWoog9zN2zQbmgRWV4lhhIvTHchLRejUX6mS4ZLFQQByJMRrLk0
2wbGBOoP16iNl4XfRRd6S07OE+BDl8b1Ld9ETsDiAX0OQrA/sYs7i4z0N2Qm0V6yHe/YUJs8EKms
Uc2yEYGV9KO7/lS3q5hZkbiKbhCacOt19ij2e8H9irqnBw/fLnekcwEeJRR7OAcQdTJ12+fAW27I
21tf7iG6DEg1wnZepTskBMVLlRrj/QPTGr2JZU2RvwgIvbKw6hX3zw3e7NFcp2jKX+97SmJdYjXL
zutBp6VKANHvqA664urtRGNeJCI4ldR/uy/4nabMj6P8I8nbExHa99bvbDVktFJ1OZXiFjhkCnhr
bMO+yWeAhGkROj4bgBoYr4uvtWzisxISgsGl2CY+5Eq7fHISrE2bIOdinJku8wCzAhA+xTbv80P8
bRzCRenh35alJqAiyOKEQLvfO9oHJyxGLnrPblAcYkGLQbqr87Ryeom45wC7a6xgMNbYtmH221nK
8Bv9iUB+Z5C/5fIpBWBs9Zuv1pOm8yFKL4gDf56u2jU/I4Q4Keef6U/KD/71Q8vgQKa7KYOYKzdT
uhdkDBNPG+FZ582ljslLC/N+N8/Xw/6yn9Nj0DaDiEwI7jczoMUvX7DDy5XkNRcltwI6LGHs43hy
wTIipYKs4wYPZLglUDyjtS0g9x8piMLM6CQgzy9Wc907MNCTDQh6SD1gBklFdVnlDL90NE1mfqFH
bmO/KkSDkI2nkKepuWUG0H7trlVOd0aDZ+A1DJUoAdkvWaH+i3feGejHtCa5ZbO1qeSAdIGuhGs0
+9WOKlWa2JDOwd1YFywp58f7/NuE51SEL6Lg/U3MHmssnU34JdudSFywLslUXIU/0RtPytC85hxP
CMd6cJH0656wzKsYfSV7y6EFDuFBrx1xkyzUFHNg1iuGbTiGets6mDN3L0KueRUiWnY3LbEQzMxk
TvaJndw8VGXIyPWLugVM4YK9xQCLgs+jR8jTmU3XI4AhJODHOpdvU2YYdkKAxad4O6LBtwThd+Pw
JCqXwglFhuh5USfhnElEsJrt/W9o5oYi1/jNFUx3Tfc2PJlmZnfMeEUIV7RAwhtF/sMhTO1QzjuI
C00dBWN6RdpxgMF+WfOeob2RUdBq1mpgBkAE92GZjCgp/1iYnCLW/rFJghAEITQ4mfks98/mj0Bw
iHum2QloQjJ+1WTX2yqNRJUyiTNdCHoXIwTFG87hg48LH3FYAMvSHKVYOIxaCTPjUm0XFz993uD1
GlWCM/1lShbJuZHulpZHsPTWEhSv7zvFVXu3rODCaKxvnfBtLufMu89jC7nc4Bfl5uGZglH1gf+V
h+WuFzRN9+4R3MjtzZwehD8Scm7KPnmGzifUdpiPs5t+ZiDuThwsju7RUoKGMyjGAgJTJNMYTMRG
fj2Pa9ZHjF+/m98d6cOcssF1DrnlyoAHtZJQFjmMtwQOOiDrvgCn2m8OJEnsmvspH+6POM816ksE
EX7TuyUziV01N9AXwQuAlDXvb2pfNWapp8+sX3A0+y/HcbjWAoA+ssQnl8LwQweyBWCkAabhjrz3
JLxd8C807V42vih8qA/oPBjDEm5wxm66PushuOZ7iHVJJUAgerzUY37KntW6dr3ir0oLYfV8Kufk
sQ8E2LneF4+FlnYUfN7eSf2z/r7EnNShAPvjd+GXwsCPqyRaYOfpJBUoMlqdPbjLTx3bk1dZlZqc
Vwd8ICn2WUL69MjJz2Gp8EHI4HP2Gd9BoXPPMjrJh0CsOUxvv1/sP/RslWoj+fPLRyKGa2YW/nW4
I7aF/UxkA4zB6SBGsUQzYczfLBiETeDkiiwv4Z7oSg1pi/ca/aBSVl0vYYhAwtvSK7d7ooziF/Y3
J+IMpfwsKyX1HNlM/3RtzCZ2sA2gG5iUJhKlnV+AdTXD74cjEpUsRIuIUmgpJrGC5LQZjE1y1zS2
q4FgFBAtZpN1oPzx6szFpYPGcE6cegtaYA/6sG0gDeK3s6Ysa1icUBOa17nFA11Fb1QyUn3QqX9W
ySJUn3W3j9GOEEWPXJtLLk+CZ9XxwXZlitPEQYt1+KwNQ77ipLyEs2fF+W/Og1I0oKquvnO8tx5e
cBrJoK7RMhj/2okHmQNB3n1upQ9YIswNSTj2SX5j8TReOjoGbewHY4HwxKipzQH6VJF8Giq0tf4T
pr5dXYdmZrAsApqzjcbra9kVy0OOpqOZpB01joHWkgzeTLfoaZe2RAxYA9+09422dujweExGtoh1
6PjqRtGEhFCkxpRn3of3tegPl8/9AMS7+guaJZeEKud0047dTRnuUHbKWx5I+CZSBkqZZ70c2YUn
ZwGyXvQYBWcwvPczdGm778XdSOzeHq33lXfXOOkaY3j89gLrVCbTzvvFWG10e3dbRaqLrdEMTKX5
0ciwGrQd5oeXtQWSv28Hts0/cPR4U2vBeHWa5DwgodRQPtN9IswnClg4rvHQePzzaAYV4I+8TH8B
VXN0RJ9ald2Hdh1p5jyB2I+fRs5VTC4Fm/WiyGxDEbaZYCjg/mAjddj8CysvxJpnMId82VS8a6m8
/suCdbq8mDlCj25BdGCZ7nw410QJEdsVM697I3P/Ndbw9gFLOjfni8H6ka9Wdd8/mv2hDaiTu9l1
jIxxeocD6waCiNmpNXPzU2SZUELGYLhUg4UE2+E3udJ5N4Hr97qPn0iYXrbVhx7Q7q95MnSC5uEY
bBl8K4DSlClGAKtYSCST3DM9yIsnI4EAaoriWAKTlqTuEB1fXoaIJosZTRd8A7GAhvj91j100ixd
BCngNo5tmD6Q2ScbQm6BtysDcCQYvxDT7oYsJff/fKwCC5JO2puu1Oc8b1U45s8QweoQ7zrjGYmx
PefNr2NHTh2ODGRMtbjZO19Ktm/ybELFg138FlTPDTtE9OIpSYmdHSeyvLPgZ5SC8VdljRgfp0BW
GwVPa4Ghs+dHeV98adKwc/PuML00RQ/1qhAnNfm+0XEzv4Vp6GdeNUFwV9kBJWaDylmxVSaL+n8K
txGL7kQIL22MGxH4NsIjDudzFXTNzlF1vuEMfMV01AtfkQUs3Nfy/MMrWgzZT1p1xMhA4qGjQqmZ
RGKesDxfyJK+LYRs4vZUlRl0PkqexGVDreFoxn0mSLI8Kxp82o6k8MrdESLmfosTTT9JcepJUnwV
2D/9Iq45AW9Sclzu6azyke1UYEJvR5ran/uLu3yC/3aiX3ZIR1GwuB1g/x8NtE1Rc8+NWCEN5Yxi
0qHpiXWYlHIWDOeeb55Xkv2G+BmM/GvGh4pom2gAILqQPjcMWHYsa2NUi/+2d7gd1O3ezabCr9Ej
TmILvGhPyxUudh7lCKHCUAK58wBAe9Hzu7VTne0SrU8+sGsAry9oYFZ/kyNYdsOE1dGHUMQSnZjj
HklpywZfAC1Y2vptd7GrhIed6HCtgQXUQRekRSiidblgMWokBrcHebSwixY1+Pu/08ThsE0MgYuY
U0whSdTANu+8ri/vwxzt/2dUSxc7YETRKT2Qna9vkbST/Vq4cfNGmAXAQTUn0UCjM4JjclWRROVp
k8C+rm29K1g+eylq1xsp53f3cQnO8f6qkXSrpEbFKYIU2burDZHEyz0nD5oUve5xS5GtAW+fQ3Mu
d/wAxM73o28zkZLJ+Mi88ZL9G+kGKkAzxShTQxl3HevGbOpVI5ZAgR6gMbOHXuTWG8qScM4IjNpw
wMe2sj/d9UScsqzcoD/ZrTzmoGGA85VR4ZoVuvGVn/cQU3XXR0AWP+scVsZFY4+6CxeA14n3mMEp
AJJ4KuPHA6csy3mHnEhILzARJxD1BS1TuGwrSwbZbMzi1e+unOo2nvpIfPxd+BzmIp9tT8KgKVC4
jejjZWO6FNRAkFeoWHgX8w9oLF+9YLXDCYA34xH7nvhHyt0S5K4odscPxI2WdgaxcUWYlLPtCpyI
ZXvyDnm5dH7froqqsUUXTa5p5tj31mr472ODg1hdJjdaymWGVRz1jC6B1ApSTRHm333euQCcM7v0
MyZT1ZcRotZ+uXhtgnqFL1Do6hTtjcZONv1GHROvEcSopBgz8UXA7p/Xpu/6DKI9xhvhnvrejWQu
QCUG4AUZKg+EJbbcWvxDYBwfFc1YxW0f7wF2Oy8w3Ivuy7mqUiTNLTzbKQHKPU7MY2d+z8tzclct
MorAMuyKK6N5PCxV887Le/iN8YgS7OSnHu9D3hcNiVCBN4EKTxv1aw3SIBt2tx+WuMjI5phYHQeO
fpuh3wwZh2Cz4SJyDVjA3l8TjY1WFUCs8aTagcW9yPoHmCo77QjKwID+NgjMjOTM/o3VIVHQfhLl
y1iYMw8PKotl1hNq5R0JKc5yN1or5fl469Y6G/XkzkZgrcyDd96bhjmZ8tQ8eo5UrH5A3/K7sdZa
8LANq22YRrIjQ8vBOcd/KeZZG7ouP3yHVxkEhbWUPcUHSrwEDzpbx/GrZrARsnS13vbYqC6IlOKQ
w9K+I1x7Zqc25l4umLUjTPHMh+UJp4abw3wLe1yUEjsjPgDp4OtmUc2DqBFCWednB8vWfUVA0jq6
+sdTySp3KWz5R/uTcS8VVIbDH8rGb0QmsaNbEcJ6fEkcB+76cgJczBOfrLdgRecSgfxPK9PveiFH
8fjQ5ZwQ4uZ8+7ZqdlgDpFnoqfCf/i/dygDCyp1qkYd67nPzBXCIrRsoh74yL/NmJeBTRZie3psd
t5qR9poFMv0yTCkGz8TlzM9qxa7p07DXj4I5d56EqY1TIRGAt5skF8klhCdSqPsFgEfeQwmwVIm7
8QIGonKCz3p8pptAI13mGf5Lfe6L8UEg4l9fDmqiQOCP1SlBZBqDtFAOoo2J3ei/JGyQ74gXAs5M
P/tRaOD0K8hVwfxd3/T/pX4jheSuA71oehk3VoI04tlVm3ZYUTfUOD5xrkWfkl35Q+KLfxbMfFDJ
EB2tyw813Fw7RqY+9/HJVccC2fOD513NdStzrtXN0XwpngGwtrrJTRWank91eBs5pC3ry6H2XWqc
cm2qOLM1W0bCIm0RaLiBNLklYKX/Mn7QnevQhCkiqNrwxJCfmB/ATl0+Wbot3/RFRSsCD9dF3YTt
RDBtOe0+P6ZIGYCeTDGuxgl6noDn11dqoYZRUrNW9ODkBMi21YqVThY26OJrcS6x5TMgQ8mynr4s
o8f0Ps5CEIXVz5vk2h+w7f7QLmcNWyVPp307ctkC7I5Pp7pOcs1tNWpyLJZyNaUeuyeiIkzeVirI
Ne8yrZmbxBoAHONRtunSMXjMC+7auBsMjpqHGZibg1M/xmzRMSrj5b/Q1jwGPJpVzfdHlizMUjDv
NlsXF0HWwEIv/A7Ifqg0mQZV8iaS/1GwOFu66pdAPrxvkqMscJMEyYz5xoTmwJirVYQZz3GTNXo9
TYH/k3VAzuu58olYyOQc+5BzRdFk/OYU960YF49J08KLOT1rsKdG1g9QXOVhxYLsGk4i7oysxQp8
rXeNPb5yiOQS4enoLdQUA3tGJA2retlIrW6eYBOzY50OlD66T5tvhvFu0E2T2HjuZYM7+KF6PGWS
H2ngC7ZUxCciFVJ+RI9DHGFoHAgrslMsmogbG+RiCayh+uAb8bDlhGvkfvEJYqGYsqDBAX3kOVro
RtEDyLbFCkqJlxjVPD5dwu5NPsxzo8jg9HG69yC06Wpg2Ct04LP2YhuNSZ+j+uaOShZZawkHSCA9
M30egl0DmvvUF8THrI6HpBRuIpIdJahXGYBOj1rChyhG7snTrnankVBtgpaEqYJmOiMhT1j8iX2N
u+8v/DVaakFr2uPn/DPh2OXgoN92+gBqBDuUnCRVSGUeIFFILE6n8kaANdDEUI4g8WJWZQcxI3nH
rFQmVHOmfZy4QGcb3UhMNlo7DM8YBasmCGD0hlh14NBNG5ys2bzyEdgqpElu2dCuE1lEQz4BBIIY
GlVObsqqIkJNuonO8cxQ9v/HTosWTwgPFlFZOoQsGh8ehkr9gK//2IPX4/lUTWbfxtniRX99kfHl
00UO7RbuE0qNkWXMJ4zubpmtZWbLWsKu/VLaHeUtBHhJIhOrS7e6FzD704rC+YUPrNKAaE1qz2UL
TpTw3a6Rco9+i6x5KVpxn821DEfFDy0PhfkRN1/W8NItPTyFNSPqvakWehugKsWTort5CWkeNfej
IY4KUCSNCrHifxalVqXTdwJLCXk41jdw/cAlAg1wsWH8j5gwWu/IEAU2EGpkKPJDX888DGVrJiV0
+31LrKE8vPLtPSwgg1KoWZzcprklVbjqCWYfrClkOCC1qgWKofCQZWnorn+fBbPueUkeifPHPVge
SSvXvDnCe5aycKd2AGJL/PPvElRExyq1z9mQ7yrxd7d77uaF0hGSRmf4OLriKSzaSPr9MA8LiUn5
NMecLi6gMJqMuScASYy+0nHwP28YkUXPh+YFEjo0JdIO/MIjc8eAFFIcIVqZ13JdCGlO1apTlJhp
9mzKEtHUnuUXWmjYhz1bsTyC51wfNrrf5hGwdDb7yEeU3xINVGQ4I2ArBHlHDgKZwgJ1QAAexYzr
9q4xxDme53y1fBnBsMosvWU6VjAWMRzWKJ6SNJflEph/EuJaZVGM8PP23B9d0hdaUSPCVq88Cvpf
jYa1MUJIHCLXmNm3+Z7RBtcD8VT4BMwXZomeNFeLCWeqfuRULAOqRXyqQffJclhZ6W7M5lLqAt1U
bOHeZytjwJXkYxYyXYYgmCFJNjjlOQfOdDaaVy0ogVrNEkxECvK6/FWvwf3PXeW1GP33TrvfeqT/
nquMcSY+P2b/BR5gVXiqLR5iyI09HqVa82iv/feQiYdcwwn667pnfMd0KPdbkKCCiBFfjcPZDmw8
EdgxyXkRbo4hfGT0yEKmhIwBLG30QDPEkrsBZSL4EtLYx/Zl362gG0Og151Z4GS7zdYZP8ElWo4/
1lmxC2Wqn3gYb3dFLWTZZHJ2dBh+8MzslPIzwJISntgoHZh7dzcZ+u7HzFGNrjW/N31aeXYrFer+
EFiXnCa/uJReMdUwUHhpBrx7Cxm7pq4uXjhW5sT3mpdc4xMlU6obqii0n/EXn6/o7o3kiHtWkRWB
H9jWDjbPzEEYIpJK8GjOT+44+Kk/DPw9L86Lg58YOxxFyRuFOjrfJcK2vOXqIMaF6tLKCdvcg3Lo
mTHOLi1UI99fhsANXMv6JXnCy13FX1gvRFP8qbTYuacdZoRI6MygzgWFkuAFmNgBixck1WQQ0Kmh
KcoMckAz8aMaMQ/UYCUEfMEhBMq846wW8WI94Au0XoL+uGwZ5VOej4YMdhUq5zh7KBHm+Lq4sVf/
3mH1w/+e5HqC6/DUb8yKiyJjTUuGFJgBTWUR7Cji0bJ5mpkOgpg6rGqytKbUg8JBEBdno2R1H5XQ
xg5qocNJE+E+KD/EG7eX5MudcGjkrfYUVycO78TRIGFWg3txHx543OuWwwlQTTE1mQr5m3novg4g
7jWYYO1JqbbXMYu3gTl8GFGdVTvu7eAgfZkoUPkzO4+KtfoaZBGyUvrN6lww+K4bbZGlCK+OPMF7
DgTHGEekpkJAzt5xFDLlhcv7TbePWKWmjY9hNI6mwR0EX60Gk3lcAicNuP4KAjsbLAWvs2SG5m3b
KTBoBpkKDw6M4qHBnuTvA1KVbCV8ZmElJR3MU1zIFFADP3y9hShROFWCEI7APSnIZQv8Jbr3Jo7X
4SDq3QZNKWqLU9j+ji0rCy1SCiRCX/Y7nwptrAgx8N+pPk+LzINsg0cO9QsdXpNPtECN18PZn8y5
2bpEyk1qQ5tNDGzNQCiHMi0LJ0AyVYe6xchEawSo0O8SLAaUU17uyk1XmcKBhezCiTANtE/oT1Zt
/QEPHK0kQs2cyczmH09tWej9Fgr3XdEh9ukBZ0gC/N/1adLwh4zT9zEmWYjrdpRC4QgeWeCRsV00
swL+Z4R9Z6Cr0rv/Ix7LFkg71tt08Jp38jDq295leUgvO5yYlqqz15w7Cxah2Kufd2802WkRM1RY
5/PpDmyrVsGa9Vr6CndacNaH0RfY0S3UVqDaaz6r12Pd+BGy2HHJybPdRbzaYfJD/YaFaN7Ex8PM
DyDQ7stHeCX+ZhEzHgylUnQ1N2xjjeKZbxDqKSNvsigAuWqeSSxgnCZi2RjVxbn+W/LOs8LsgFhb
civeb/TAhbyrPtLpQqZYeOlcZ6YFMhVLUXhLREnHckZnMNNRO4S6ECydAF/J0kNMmP9QjFM1tORA
a29ALeM69DqrpVwTLqPIjLCP62qZxm6AcU82BigSvaRuwGH2ISvR5Bw4Pk8EPq0c+qxkVsrMKFPC
TsbH0t+QfVXs1DI0NsYtcdQrO71UHqQWvRUAKTCXltgJu/joiXbinC21p3ZPkPgs4J0SF3B7aClr
9d8+0lALWDMhmX0QPOUmq9MFVN6gO7mMsf3kiw5xwywNWHPpaNr1+5i/4aR9dsfjspA/yvafeFAn
ZRbrdtMDhkofFL0oFYHHPsp0pCNTQdBwVRvkgrhhbGknYEujqbvuwK5VqS8SQ6tfKq7RkS9c/onh
7XOr+Fr3K5aYbHirj8sZydIO8xG8YUrZqktlQ7Jlq8xnwLAXna+SUmerrbmycsWQPEdS4ugI27z5
D5V1Qd/CxmhsCRGRFrPQpOfW+imWCZzLSlM8vM2v+LNGjA/7Q5VzEpnryyZCwrTHi9GDRB3MsS4c
Ap1Pbiz45PajhO64bLJWJ4aDoYxTQTYKu7ngRQ8mxcjXpN6OMIP85JG42C34OQYQjTsIOCTU+zXB
l9kDbgYoYwkEJQlUQdac7xbp3dd5Q112hSOubGKoBEs7Vv64bNAqDVUn+ntWnqMAo0RLQDYqNyT6
Fig6B/PNpcey/S4eEkHDtqntiKu5E00Q3AnTOLb9YgLnwSrPm3kOqATXqIquWxPwbMAhaUW8bZlA
kEQnb+RPFRoWeLQ2M2Uh1a10keiMMLjz2ME3wT2VRe72c1telrBJkZVbaC/hnffrAFcPrzbgZ1bN
/mJJjEUwCoWXH+iTAG9BfCsw4kO94qOfREJpO85vgoHX/A25fSqxtTlsTVVydbS12RtZ9ZELn87n
NNR7f3xHnZLp0pvw2hBPV43gOXYvRygrHIJicqka2MBXgTwWEzvtE5cY2EJit0L2QLlUjlBmbDc0
6ejBqwmq4IdXf6ruxNBcT7C0JDOGqHWjKna8UkDxbxL13Jmzx1LQSIXk6EbI9xVZAa8u0/zLgpjk
ktRKwNeqRCnKp45c7RySEAfH0BZ1aEhDoliGo5Jys7/+cf4akDfHCX8DGO41YfEjxqSSSDZQPhWc
nYF3FJhWptbf/mqhBadgzzO+BJ9jHpP84PAlE/aWUV4cN6+jJbqpNYVMhtKPQk4AhtHE7ZrYCL7J
WswK5vc37N3GLvncFrjr5Indi6GFqZEUApkkOLIC0QchSRS1EZl5tru4SR1gzMpDjBzyTFi+QpiK
p+r+WQnHTtf3R5OgQyUgql2Sb1KsEZnmR7CC0JM09HhReChaxnlDtWVp1nBbd0J+Q34gzwf+US4o
BPamNi15wqtQo53F74JuxvgXwRei6DNSVZCkXiHb4wJuaqlUHEk89B/s8U1ufk3etFNTyI8122Uy
i5gNh67gIPH9ihYofaFc2rnfMMBEXs0ZJ54Gd+9Cm/0ChJkXTXlXzRQp2FOs0D1Qu5Rma6NAVMwY
pYyLIH5HXXqbXI7+57qtRtS8OjNsvE2cB2vzP0u8RCqPLLU0O/4mmj6xLe6XldqmV8aHRvqoH+B8
D5va9FrZQh5FWxQSsK1AeL4vNWvbnF0XYcma5fELvbRuZdvW56jxvTfvIVKmErtzyXCKKWu5nHgX
qvPtrba10goY4CBxvFlze8hANsVXvpcMjoH1oKxFiwn7+80Jmie694ibkv+FoEeW5yqMfiALQx3A
u3qd8M5H0P4WWtNW/ReFkcwWbqrmToL/2C+z1v/Su7P1whjKwCaXLg7iqmT52Osjt+b/AygLbJQD
Dpq6j4Yd/WnyX5m6Z6gHJhV4xqsL7+qkND6MjvIBV7DEj8gZrBtxCD1tehsXlaoXYhgZ5Pntxc6k
kI18KtAFhH99FXdLbyuco9C/WYtHgfqk/i7Do82Hu4k/8BKIgroM98M0WDvXFpn8T3B1KbUJSMPq
dN/IMANTyioPHf1c+m7lP6w7QezqkBW7/IUKn/ZqyoKzAZJhakyC0lsNKr70Fiew/2a+8ZVa6r04
emeLO8VwkkJsLvBUiEzY3s0Ag4fms4FMYwKDLPvqFyyGX0fFa8XDkPK5hm8PgArBFar5jPbefTLB
Es0xTbKwqQEo8wmJ1w8NzOzjazdZ5q4HkEJOdX9QwjKVuvyzpYgupRAbEDCwHD8f2Z7X+CDgAPS2
oSxh+zYnLQJu2LPiYxKCsYyekXtpg16QVmOcdwWaYCuXMF9ozYwVJG4UNMGJS90xogvbUcrpuI7y
Sf1FxIpZwBHDBUrourNVIIeiuRCdHoyQ1elvTOfQGi8ykCRi5lvadzqqvuCIUCxogSllHKN1dR5Z
tIycrj1cqj2gucVKbKhQo0UzotoB/FRPungQjG4ZtdjxeLYiUTKwodELcHRj68ufSOIxwcEd454o
vP2I0ijoyF2Xc0pf5B+JDTJ2RDqh+93pKbTtLwCl3WmckEXrLFu7ukUwtnRfsrrL1mTo/dVIB9+N
I55EPKQPOA186BxVDn25gKKe9KlKE7g8SRJRC4P2zBzYhGbaVDth+/jCEgpg/RIqXZQOwmSLDagy
zJiHuoR2S23ITsb7kj2W2tOxafHGwbsTfy4E1EkHbspx45fCaJ8gEBtRQHwO6zIPSjY3T6GYJAGP
Ps5tsD1wa2rJeTmHgpxkr9K70YAOFch3x2JsvoUBah2nP5sgrZBpqKs4CwE+2JP7aw+uWYhX39Lc
NwsDXxhVl5bbQlVhs7vHtsyq0rGczETnar3CujVfhgyuLtGCcajQQvtCVrwsDAqjaQ6AGg6Z4luN
gjAQ+L2C8tje7XTTV951t6eoPBIOEjnGA51MT7+3x2Ce4SA74YmB7v1Snu7GiU1g09eQopBqm9zO
IPXHGwu/mei1E+MoL4JG69TNyR4BiYK/PkEeIAbJl8IcCDJMAND7TzLsbrfQAiGs5/pUdMo3FIvS
8/iFrv5kvz8lefsFx9zy9iBPD1Q11GkVs8RIJVzAxFkLvYGz+CxSmYy5AkcrGlMMlDFcYjGz8QsG
rmiS3bebRs5JGbuz9ncCZ1z5LCpfVB6slwgcYLnj8wWMI6GqfzmMGmnfurEfSednLwbk1p0HONRg
0HgSommGx0QzU8uDDyYquQPMa06Sj/xXXMO5SwgLJFNR+WKz4wgMap0DjoWCZN1gmU0GgDJPW7EL
HaBl1QQepZ4QxZ0Peyd09XOUFUbNcQKTQ0rGOlJCefDLxjzvfD+dHRiyATlQWywhV4o/i+C+ejpF
WVk+J1NBKF6YIt/zpiaMKq8x+6yZ/236s/H+CWLeu8pBV32tQvA+pHcM2zGqM0IYpPp8Z6ghz0EF
Nhq9IxYwDNhvn+KS9MjgiCMHus57DAe9mXRFx7MnEHX42mGiTnmGesK3o7b1D7J9XLWiZjDCrP1r
pUpYhw+4CbCjuztapOc+F1CjG9hud53vCJVZJYepU1spsbusyZC+DVqgVXxxz3zXkwoWzei8lITr
c5LDN8kds7UvwKKZYZmCAdibHfpIAnAYeRGg16F3AxpLXjpKq2qEosV2XxP5YKtoepKc1JYpZIk+
RTPDcbcJETxLj6IER1vPwinjRxNP9mUDMUWBwg27LkCSbxpRWgpaPis9326gVQG3bMGa+c8JzzXv
1xXxUky83Y5K4ddqnFu/tYK0rpjEviX/8wMF6/Rm/bm5w0fLiMkErCgocPc1HLdcnDzLODTv07Jc
LUahIfPdSRYwclzEXatYr+jY0w5/8cX44ApJogrRnFBNw74e2QLuMdy/ydPPP7jmHofq6EuukOmB
evfmgyk7hWZOFaZyr8sFLAwQoxrmgpEzOYJeywmsu9S5Hpro864dvQZUkLrZVtYoFAHpy5P2nAzR
J6HKm4/Jf5R6jTtYa6/X1nYXAqY1kr3wH3hTUBRiuADTWZ556EQEqPBEk0Xc81GSbe20XcL1ymIY
0HVIJqcsvS0vy94OVLQHdIDTCB1xP3drRTkwmg0PkojfthpN+rdtnXmhU0vvdvRKf2SkCuX88VaV
4BPfBqM+3f4S0LxupWZjLuGidH553o9YRwSJ2IH4qpu5bl/HYIxpw+Eldd0tEXdgwk1rNwznklLg
6WPVze+CFl0tKya08uu93zm6sf925tsSeMg4HKGR4E6SuYk7BlOFITwHPnrhQLOzaNAE7kMEfbM+
eUG4j1CHCwoY2/cMVbTlBTIXEbyc5sKGb7t5CVErSXfjEI2gR+54tuyIjTq9qXsLOx5vTH2W2m94
oXtL6b9WNyan0HBciIrfCGR7ZHKGbMKDYmXhqTVvoHbX/vVXxIOhxalbWnTHXQ7qteUs9Hu7psuN
p980USKlxGJyQ3tI9qPmpR4Ul+vmjpTJn/BKxYWQKO80rG8p9sYNsd1fTMV0mHa1hHNiySLTeGEs
bDiU9U3/5DwlmViMYiFKl28HE3AdwLDDv/BxNNd9bvHRdXuIcHPQRyyzXT1KaY35BBFeS8np/krD
uV/uI10iRH/tuNchixFnRhuQdIa2pNyTAhnlYzNKJdjMVpbcKGymyBFuMZO2gVmscUeubKqUHSv3
RCxQZXjGOIM8dtRRO9ujCqn9qaXAmQDD7y1Nr/Kaav9MkKyWCziS7DOKzJJy8LFThVqTMbpxhuBX
8puNxXefKFVb/KDPwmwsPaNBNq/8Tv+rDjU1RFNY7HXQXzsCSyR1djRc6uTWMm5+343GFB2q7yep
BdRY33SQs/ltbB4G5jPcP5rMCjutY5Ipk4lpVW9fU9xXx+M93ufJKW6g7aYmohlMsFjNRMrzcFij
IJw0P1OEAqJ/ex9s2VH0W1uAkCu4YutLw9RfZwynXCrpt+cjjLZbYKQsvz2yHD0TzJKQQkzFRKal
WkUe4AQxDfRFhsS1fVU5oduOvULq5KbHLhOsJF8fk7WWKee7b/kYHu+di5zwHo98UZJdUFniP++8
nV0hde218tAsoAgLcIsji5BO0bf+u9f9DJGI0lG16JAzAOxw6GlA0FB4OIc9KKKt02ga3JtHsg9W
hxutFMPCmyh4MAoYPS0FGh7Mu2xFon5h14dAAGdhVbHhY+Y9RJkkz5tR7/TwuRMLaWWMVN+8lfb6
FZ5E5MQeQb9CdRRzh30rtSLwXw510T5oMPSoJA9mOtp7kG7SbV0ljOKiMIqdVnY+i5VOajjlqRJx
mFmRZ3N1NPZOHulxeID9SeN+i5QOLqoXCBBBC0Yp37sKcCviHSWEFvKyxP0qWjllmw3KDEais74T
dWrPEUjNjInRkXuuGvM0X2tBpNZhQtGgyoKbT7k0VQiBuTo7i1zcvv+ri2KnRNhbHQFuNCfXV8n6
g6ROJCGVKsAhnMTK0XDulNniEVldJEWz+q+9nBaCBKpOdaifPKfYcaKfqVimxm0RTMyQOWIBXBk5
Ci/wCm9AKj2DAPoUmlDbyKNx0KDZHzi505/sBJ8NwREgMyPwryJr3LnXqUIN2APd7J0O45k3bsOz
eivTj3KS+F/2lTAnSsuGOoQFDmMV8e+y9ZGDrKfT3a2r4tDS9l+ZmlWJpEQQvqIG+nDNiMhByaqv
guvVd+HFMZRhqY8Le49odisK/r9IeAsqiMpFzdlVrDxs9iFlYVepxJnLoMXrUfA2eKVQkyGSRwae
mATFo6DfNWMNGbWvqvI7rw/XJF7Y9wQTzfbB6E15gkVd0q22JrqPaddJOD/M2IIIPrHXeBG/k+wx
VlAV9kIDHhguHZa6BIupMjmbTAnHI51gwCJhxAX+QpoXWd3I/LVPeXa3nN/OhM3MtlNRm5IVOPFx
rw2vP1xNEpCb1bE6aoLBC0BqmUZt4cEDmIoUZ4CocF/UDBAKwTDbnTetrO9AQ/wQ/QdT5L3F17gJ
RA0331MnL5ai1Eygk8DtwZoTZz2dP83mwJufUgtc3LBOpYEsBzmweY/rGDKPIn/XwTeagdVqFMws
LCOVxB30aDqttdHVF0QGusWAw7DlFfI16mbVMkiaSPtJ0Xt85A63cwkNzflpZMfxT5Pn4r18XP1U
ulfIwl8eLyNLSZ0f7ro1PFJqCjrV7VAuN4YXHXXEonInbm4EFm3xcPgetzDjys94POMTA45jdMLq
KpxC5Xx0gj4M3IjeG2Nvop3mV39CgPiP25QFCCiVmHqktvO/ZSBVwMjqynQLi629LW3ERpvpo11U
nZfTc+7CH6DUcC1J927G4o7eBj3iv9V9p4WSowfPhfOZYIDAGEd6q85lAfSkqfq4iqnBPb3fFkTX
SVk63/dDndIPBJoQSdKezl3x1y5uRswsUT3JE+mVE4hxO+6sWlrQXZjbyeo3YOpiwEglK9y1fyQd
cEtPYzEm36iH53vnDCbxDff28xGPuLzIhJdM63f6EP6fhV6B+ZSSYlzt1wBDItGokGDmndjdQ+D5
5JRE4Ya1rzUz4YdOi+CbANkQKhrbPlLKa0HeRcJtldcHRq/fi40+hAOMvg873IWvJ4cLOG5UeD1k
HZBfbg/L8sSvsrye4MSfcq65JWFD5CzKuYIsc6hVbOqegIrsO9gx2dtjodXTuJuK4JOHPqEXliCy
PS9hWUf3KZWM1vnWYvNWXhRyYna00aFtdMV1AX6bZxau9+HKUuzLLIhCeh5pFiaHlmu617AyN2HY
d84dETkptD+OxvLH4CiDWw3XXpfi9hmGiqkgdxQnRC86N2dWAAoNPj4AMbd5gEQQtPT6xEYUa3GP
Jfr4eCLBMEMInlczvg+bpZ6/qz92P7v7G2nYYRDjRwm1H0IqWECrgRcqyEoZX0m/ibgM1sbVh0Ae
RZxWp6tZ974EAL6mwPCkZ3qUNW9rIGEmv3mQ3TqF3cPBgDhjjO0RsIRXYv3NJ+FRQ33hchcy86t4
u1gB1VrgT/wKKYGv72Nhjwwrok3W0XNc1lSqMUlExklRlI+KflhcVF1s/aQRhdDrHfTz++kPkA0P
btMQMXgcRg5BeLwgAdeTsX/igzS1t/snscV+U1dVx1xAl56ehYy+M0DvHnjkoZ24k/GzwcEq1xHz
iVwup4QBQ2LSlccypLNjOEZXW2pGWPGjVVcEU+PH4tp0zxMe8MpEgC83M8qnmkzYSutKGrZSbR3J
cUyCOEXuBCYzeHKw5DvHusT6Ga3wGZ1Haz3p6L6A59jcQGCGkd7lsHm/g5RbJGzEOkDKQDJew+Qx
HB4nMV4NnTOt4fODc7nBaYCV8oRyiRIH7Aeic5wGdPI7Op7mhGmiIJ25KhfSI3eE2uBGCVzTA5MO
bGIqGZybbGw45mmaapueE8nEExnny4qKHmT5IK7HTtdtrnV4C6RUtQcP6/YXhmNfrY4lewu7PmKe
+7zBlAJxbF6pwmFmdFXWck2EsrO6vHZNu0YNigonB9s6oKI79LCrFeRb+gF3AZk8JF1lNCRav8su
uYIp/2E/F9XOvnLK8zrWseuqrQRh1qDGvK97+q5N9SzOdp5BSxB9JOlQ1dLUWDap0JU6U8guk6Du
OhDae8EVDKNoT/vYCA/YL884NR6xgU//tBZOjMpNtKwGpEE6KvtPheNx8+wywctNjZKesppQwpqk
Cuay+YkiEFjnEbO2q1B5+/AFkx8OklaVh1fSDYo34oZNmh+LvyMpdYs7kiOrgYXYMQI7I4KcFrJC
GocNcFeup3L+cUFes6CYKxa74TZw1/RgXrZUlYVjFSAKxbgP6lND+ZHf786xeXI2p/Pn3nvvIRlG
nnaItEReqZnf9ie+Vu94zVDNcubCcObcydN/5eoHvQlj3/D0Ty9UAJls209NMl3fOK0k3TAfl69K
BeYnHPLJWE9MXePB1oHjgfqj8y+o1tPeYVck3OD8vEMXjIlhfdmfoHwfOwjkcC33kaOj3FQ/4nfr
W3+94ZtJS6JzHcszWv9fWDk5kGE9oR/g7efDOCzXJ4oCPhgHh8Sl/gU+nWWVG2QClsHB0pBkXYyp
aWng64y3SQw5U6kmBMQX0/OQrurm5N3/LSuizzrWJWxamz29OQDeoS658/nPIhShd8rll8xmhN2V
2lQlc6rlENzKC/VzWueWYqC6QcdCRgSGFg9pHEMhu2c12j2GJng2wJ260f1pgNPyO0pXXAqYz3Gf
Sn0g5Tt8rXwCuIoiZ0T1MrcUi08ZmtWysz5elUwhXtcPNBafHjpdEeiWT5sMK2v1G9oO/s2meHcR
ib0wNquF6TJznNrWQrR82oaGNhQZYFwAVvWvMHAh0pnuDfdXmI65mv33E0c6qD0G8yfAuurbjq7t
/Q4oUHPSBuE/cf01hnvJ358Og6104fnvVwjaICuKuwbWfRb5bQ5zZv0FLebigA0so9uJbbskkc3t
QaHKBeMM+wMxud2pxsnCKY12V5dWKJFsHp0Mb8Hs5qM/LHWDgaCNtQXWTc0yJLOMabm5upbJK60E
ThYN+hV+2GsnMgZaafGq9sc1M0G3/HkuyAJakxUzFn6JDb5HDLCMWeu1OH/zwXZ2CIC1fdCZaqir
L5H8Zt2ltI3bQZSBVOUGBxUVkAVobFkexoGA1xwWm8eG8SxdTeeUq1+BuEW51xSei589oXk2wRa9
1xKK9L/i6J1YlPXBtR3n3GJIvMSQUf8lswAxh/qceq7Hr41Zc0yZLORjEHvqn5vZx/5uuPWQOzEF
HfDVNRxxdg1lr//wWvOF4oEKN/4PxIFGBgOWWBBGAIPKFXmqiH2ELpRJzirWLi0GzgdzarnJ6kvo
5yYOPaQFldjN2ZpsXIELyS4ZRFQ1lMRx7E2JcJRg2NhWOBQ6fEHoGePF4/HOsodLcmW7WZV2b2rx
Xjz4dtlcz+O3bzaEMNWS8L6Eb3G21mq3257iRI5QOoKEiAtHtGjSIy9JaAQSWOFTkrfPIFjD0Km+
KtUcTQA27HBYFijK/1/S1rafuWhEsOhx8IpaGTY1PChhFh8HFaoCL8BIgYcQQyvxLWn14Q0tjvyb
nvd9YyorlLBXpcWxMSL7DjPfxLALZpmZW0kNnvXT/JtpypkIP1M6Hb95S7YzlfKxg0Z/CJ0ECNWK
a4iChyY2fzQ/XzvO8UR44hKgZtz/B86/bAhKYzfoDDYTmPnSqYTA0aLITE0QHcyyZ6d/3UY76rYz
AgLxaTWrG7Wz46rtWLkrlxSq/VBNKTZjUkHPQmKcdvQxN3Qa248/4RYWSYW3551i/ngOUg7NfWG6
oww/qq58HQsy4aBQj1VY9EqxcRe8V6pSj0CVBo1IIot8+xIDebQyPQpeS470Rc7gmJxGUaU2ZJVT
Prs+I6YTv53gyXDGlFCW5KKMPW+VxdVh8930gBnqYDpVSQa2tpM6ZbaedKBNMOhOM/9N+He8uzWo
FITLUCCReiIjUzk8/gnMClBq5MgvzcrL+uSyfe/Pg1Bw3AaxrIFuYDD6+JeO8S6AfSF/o4XRJzY0
cf3edrcvUrgl9EcUDHqgXSB1X7ullqg7y/mBhU2jwG9ofo4M7iVd3eYxMOg0IUmIUWbGjkDA1nYw
GDgevhqVJwnTjIyZOiprgCCd/5og8kSeFs12oWiG7f6FbJAjHkxqVYBv0RewdoPuBQjUrCZBmD++
ZOmCTSVYETI0HzLyLpPlLG7JqUJMwt+4ehFneUX/HwBgCc0NaodJES3ZdypBGMbQTIfLbkhvfYln
qVAGGCScxjaodQdUN0x7FkaVWKG3g/bixukS1IMxZS2rGqQjgf20cLkdlCglToXE1EILbGIkQefo
+dVEyR5xzF7Ax6a4Co4E9zDoHR6+ulO0pgCHvLGEDE1oQ0X1DZf+m0SH7cfDPt+s+GLCZwwdLquC
XN86NyCu6jxmQow5CNe/J4PFVg/hvJR/L8MkbNcYl3hKLO/HoCkGJwRckS1dyc4pUOF4H5DZDvNd
CmYnPrdf+CVUn9eGIdYIB3ER8FBCGzG8/cOf37XLkuz+Qyg+R/q00TpL1t/ARwNsT6UdHTUTPRPc
0naOmO7A15mm0sby8L9kthxrXWU+z5HOM9V93JoS3Dm0ljkTY/+eF71LQnTMpgK4KqqkE1/KaRQi
+ZNMBJMEIwYXrg/EMB3wa72vFUOkw6Co/cnCkZcmR0NUqNKB4HIpVojbR1AqA/JPL7VgnLEsbZmj
le9mRykeQE9edua13xl/cI9HrHOE/VuiaWkkjBddePjc/wiPc5NC+8HYfjNtdSQ6cN0UCYt+4LyZ
FZliQHmnhqJvVPHT+y9vsxpQ65tyZkQ6yY+rcsHFbdzJqk5sVpenIsfzE4/XsEY1qqz6g/Pk1NM7
9uNvro/J2MT9RI+N+DLcWeIAgoZi5drdoyXOVPTwf/GV4wP5CG/aXmcj/sW/66haYljR39kQAACz
KQ2pP9lE5N+NZMv+GvwhuNpOHtqxMsxOronyS0j52qjDDT4jDM6p6vDWVQ24wJdBuZlp3R5UzCtc
Jd/6RQgvdu4DpBEZ1cuM3DGk7p8Y267I2BptYEF7CNHLupVxtSB5Ig80DBWunP5FMFAS4NXImHaM
7KA2IhlOxsJ44eGCfoU7PrxdPAXiy4cTGSIHUbvuiUq0A/hCBb2n1+s/zN5NNtkIU2xo0BAfee+J
17KIPey4e2PAbrtsBLz03cMOvJ+DHnZ3J6RmyBpWrJFLv/K2xMRHcmX1klRqrpGUfhFwusK6MuaS
OXvCAscoHSmgboFX4fD81w4Y42Aixt93zHN9NMKOuk/GUYHgCwXCeVArtZZ2G7OQdf3naB/J77eG
6yeHJBznx+ay5iE21zrlfYMHXoCKsQxamBl4WmYGb73jekZc+Pm7SN+5TdrjIvMMH7pBIqjcHodw
pt8HJqpfV3jMnqBK+DoV0OwEHlk5rTIjfK9GvhamY4FT6mirxiuw7vwHO7RXPbwvLpeYb26XIkh/
WieZKzWfYeEgfo7MVMiMF1z6RrgXzLiLKl3O6GM7dfNm8zXJFhetRNiBhs43DfrH0QcccT8RRT0c
CO9PVvZkIInCGV/pt7OYoKqZZ/eYgPLSfYmX80C+I6nrtyOalwU+UGSAa+jmuCQbYxX4Sd0l1iVY
k2VR2dAtL25Hwx1eoTYrtl3+8v9OqACtCF/aj/yO85AgPq8DQ06gBTvW2PLUYDM5cQGNOMWj9+bx
9WWV2gXpAFRyhfKiM9ms5sve1YBzKIcUqyBWlNnQQIXgXTvcMEiCShVk35s/2FvFvaR524SOR4Lk
3z8OyTDD4ciTMAASTIcOU2K9wuqzpo9Uyoeo5MxFpGFz0itioHk7NUd4hQZgdwkR72nRN/HCI4/J
iV3V3euUfnijcGUTTQir/UeptxxioFxEmDGU8gdXSn747ePrAAFoydY4WCxiA2Ea5yQ4EriBTtWn
tZ2HkqfAZLhigQ7x91cJ3FE7i0abNQUpNsU42CBx3nH2/kY9yjKTFz0CDGokPyYtLtRqNmflZYRm
pgZMMTYOPqscrlHEh2xhw6PIWnuZXhA+spntlrxNMo/33ftgT1OV1C7gJHfGgnu1cmdy6/BMaudi
kKwizzdsSUqJEbLxRW1UV084cLifo5uCgdsNQnZw5udN9EOP4cX0id/uMqDCZbw2tbSRKXFB+rQ5
ALJuHkEODd6O0zXDFxcYZKFVMDUCUZ9uPF+4+EGOB6hoB3WxndbB7AMLK9rQu0OxHOGmYCjWbrHb
C/f8Y0OjGu22WaiRrjyzmn51DHm9RM7Yx1tePZPL+Bd74EaUpssICZGzuxoc3ehWaisjdhSSCxCE
vybtXDVQXwi71IXKC/Ylfvapcg133QP5JoWlJ9epH+tlKaUHAbCpui2DVNltx1l2md9UXpHoGdW5
gMj0tr5mGw9oSc1dOghTTBjB40GTCeT1gwia++LGZWwqsD80UpEo2YCA+NnS/pl7PGENc3JeDmNE
Qkk8mbYy0OUG8agID4QCZLmyXeVBxZYdfUy2p7xgB62+I4m3Q2R8d7iUHoH7KQsKxoxwf2+F7NNm
3Lxsa0U0sh7EnheoqHHa8RyT7TDMJgq1+TMWoko7D0a+Iw2cy7qJiaw96Qcdw1a/cCRCn4izNN1x
D/jywxf7cXYqSfe9A21PGwAnfytwfSYKcnxG4mflpLWo13RjWNkl4CKOnWFn8RVQOpiXEDJkzH+u
bEbVwuNpDzFr7youoiMPm/vo7LlHCEU7bysJglO5UPI+B9mHBT+sHG/E8TUE2LJQoarAo8+/DnzL
Vkc/dqWDRm+V9vEkce07GCE8iFjY0zGQO+Tb9OEalprW2YtET/mYrfb8jRhTNba/1JbfhheiuAOf
kd0wNigAFb2kGfP52pGA6ojGa54h5vr1ynThvsfYjo91LdHeBNImpF+d0hywMLL5JmlirJfiZ+Ql
vCUbO99fabwMOCSoLGjPF5NXfO4y5QLu6LuJWnTG1fDkXM5DvQLe3hX++Xp4Q9LqTJY8/umq09TQ
eUIyMd4THevhSLOnT5sn962Qrws2uveUGMGn3qKDeJmwOrwrU+cF04bALLcla/8v1wAjKa/GeOvV
oPHiOuIejwUIa78t2QGBs/1glShXSG/noaHIWjL+NDV8Qzme0an6sau4tofxN2DjqlvoGYafhE6q
afU8g6eQTBiZ4J3g2AUjPyylL6bhG8cNYL3wX5B41RES/i0Z3AZRLSkM0BFMu/QsKo8yts7uPU8p
Y62VKgMz7x38VZWibaZxgdFb0MEYxHoRacTPXPZRuKKFLEMJNaU1BzJ5F3QacdNWYykjGzb/mL41
PZJRsy43H71cF7m/B/+Y034zIPNt2FiH209eH/jwgRz4Z7tHYZfyBx91wh8v9FLhs3/V01HMXPYP
jMVLxjKf/IbhURxqT4/msr04C2gpv6OYOankFGo6GnXggwotf2Ezl5ty4ClG1bMQtc+tHeONHMwk
AoyoG9NTzLRZsBqyKenARfZ9bu1pLTSbQtXV2wckkhd0ms+7iOxPoP/E++NoNI1ELhyo1Wr8gv0R
wlySgEXJaylz06qgKEF08ltpqAS1xn6qWe0J8d+VVIny9ljr+PDZc8wR91NBL0k0rWohdf6gunw2
7LNRjN19VpBNjTAT2bN14PA/mqKsxvSWoEX7jwUxF2QAcVobKmqoeLLYfmUSUnuYsNjODYATRPL2
zutWQgucACKEwMIfrFcMnTZ+g9Ut41/a/WR6Jd/O45CKx5Ela+HAXLT5PaQFQrXMkCFWUjigfLHN
E1GrFAqfvPZJDzaOLsUlSaYR7l3p6Mlx+0QIbJwznTt9ojKTeyRIGG8tVCMZSsvNTc65GBne3tC4
z0hVuavmO2IjCqljuE+Tfq+1WHhx8LdWLGmeHsz9or1AHdUKrI2lx0e/j0QsnehFRmQOVqj/vUnK
9WOtUl/7aQ6dqYU9zYCy1kkEWOzsiWiBUlNZXfsAKWKaym2VaEwMw1pmo99lPQ4YWayl2t7aWNn3
ynbUmMiCSkNIlzuVXGhicI5xWX2CP1XBe2PgzPQvYA2uj79MJrzxOE7hUw1do+f8G7CbwKPiSkzM
PP7yZvDh92DePlHzgZWkyymT/tO0pDowNrBfhY+tdcVfTM1ylawl8IJ584/eomebVjbA8xG+2QwS
+3HWfbMEFrbvOYHX9sKn9wG1hJjxUhU6yHKdV4n0u2L/bye4A8G8VMHKWHTauJpNeaCaq6UVbpYT
yl86GW1kUXqQYTBw0r6hRajDwW9u+Iaq9Ux8jMO+5AMcPLvI+RWiaMjGkQIzXG1+9h3z+roaBUGI
RCCVQjUbEnfg5Od8pkA2QU5GlHnrbo4zTtQ8KgSov4L6dheg4g6ipIC9HhOqJL+s0r/VDTCahLZF
mAZERYfcG9g+8XmreGlp2pj6cpIuznJSyIEakxahANaktooZDSeSW/BcRnne4tEV7gA12lRhQwOt
HB3QV2szfEgtZ7tEK80qzLgIsQpbXOG5Dm36i/nlUbcy7HeanAGAjM3cDBkdY9BlVYK8xAOP2fFV
Ke3+wzftMhXeVdB7uXEMWdTUEkiV67MT8mtNvJ41icrozY3JmcXjPv5DMqdlYl47rfVi2VuO+jch
YERD3RajTctqA6hGHRHoMz2RrPbXgTw2IDp0Ne5Vk2u4KvtbhpsnBDYU/lj4h7G8p+Scdq9bSnjJ
N0ab4hqGYVqn1nnq+wCKhbP5j14QcuQoKc8nOr70v7zEJZYaNXw0JwaE3lORZVvsV/3VbTt1uGhx
mjU7O1Tt0KK8OACcAcFkwWiXqoQOz7cGZAWi5pZ0Cd5VWQHSFEg3U6laJs7HPkgjLwPXmlIuN66J
/KqMZuX79dIGcrS8NHu4kdayvaylRcqnn8PdbBjXVYHPuII7zUhp5c9AjcZcvbiBuSPl5L7gF3Gz
7UlXc2mjZTgyHM5TpsF2kusYKX1Ofsic5g6+lB46AbwUcrmANqMfwxsWTVHHw3qnvN5gneCdyBKO
Ro1orOKWR5sOUNGr8gV6ewaM9p+UoZcFxB5J7PlEC8nOMRYG5sdTnUmpnfZRddUW1VzlHAdG1+uu
7QB7EO4Kam3Jm7/TrxwXHLIH1YSOFM7jfnee/hGsIcVtlgmVQsHAql88rgTQxVybwDB+r0MnDEpP
5hy0EKgfISQjoWTcoMbfYd7acrTPbcqAGDd1U8JePJcDhOP0hGoBJNU/eUwrncQjSPiOpjWYNril
JP3KtkR/U6fL48S4F4eSKJki2ntgT6+EsXJKOA5kIL9sImuJhZK1H7hobmRPfZ0BSOnfKq9lS3FT
ZRvyAwxtn/iNQaQhYrnasCbc6lViPs15SrbF6JUSPJBSSO8JbRERAUN7UD3tQ1i0NCVWZP3DkT4B
cmv5MKFP31gCXvuD47AKklK+5KraqPD+ei1dxCPQA+V0YTBjodEqUu7mrbkFMk+ofsgLMcWDjz8b
XzOH6NPmKS2btVkJjb1YYJFnyRsERE6/hy5+PyRaHswX3XNcROk4Zv4ofmwXfF3xF0CUZHtFOtix
5Akj29MQjQujUsEmQ0vmSGgk1sNQNfdE7IKXnf06AQ/1uV05HKrgfEtPiDJZJS3qZaXKmAYHr4BP
9FBqHrbuFo1jqN+aY0nqGQ8BTP1IF/CwdijadS3DOMdcE00MpwKWxbR7Qk/beimdCFi+/rRxbtAz
MWXWnMNc3bIfraG5NAD27KNLrychA93ypxmiJzTGqyQW+XHwOtF7Y4owhLlKNTz6cij2C846SXfV
rg7rKDEB927aaA7aLXi3VU0YQ8LcRkxmoILSQ7dGMbs2/B/QUy8pJfSZLmj53ZfVU17szRpf2/PY
uoUskReklFaSyAwB7NY2E0S6/TCY0zQyLn1sBaQdF7AS3UBknfZ79ZhIMEuS3Dm0dRySZAZL2ybL
ELqPrVzAVPNDtOUPVINphCH73XM1WyNCvw5Oh41Zm/ljBqmHW+7s2pnc6BtvdNQPtUyAihLaqadZ
pF7jTKBf0ARPVp4YdMl1oofjswDWGiORsBALSJwuUcsNCtCm0dV+Je+ivbH5NUhDwIA3MP/OdEPj
NURAqfzJD6Iqmn/f58MXvQXp5/bv6pPo1cjiaLqQMcr2M142+vcHFvpJz2Z4zul3AnIfUFCRGT3V
of9FkiFWJBUqpn68ijvtu+XRMLVCv5xw2aj8MjEQZrjNxBzfIaBpMKMMN3WasVyiAV/w14HlbPLK
fZkmmg4OTH6o/fofhy9+B+hHOPGK14wm6bISUSaVmyS3rmdhfMX6gkS4xEk0lhf694z/PLj1AtIm
rvoemGxy0zvbOmcAa+r8mHbg79MjbtLoBs3BpkgAwUryE6fGPX13b1nD3AeUXKg83oJpKEw/qFgf
tGOBmeF7zjx+x9sT3ahbzKXOo0LcvW4Rrw90HqOnj8SxH7wgX/tPUlcIQA93v4x7Ses8DvJQmYmV
zu8pWuCWu0MonimGXlWji+5usmQMbm/S9UzvA9TxrTLTohkpBt4Rm26YkOyC3GtJVCUtswrE1mPD
RyJ7jiLQJO32bv9atblOyKFtQRFCsblVp3hpsVeO1T9k9F2Vhe0vvgkXU44c9uOkz+cdqVJgqqZn
7Jw7G0JusFWa0GeT9p8DQteQyV2xQhfyQDKi54hpXue+rYufW5N7KpufWjKMLCJNdMWCJ9+cxSRl
/KGxFRFLWekmflz+a6m4U8S8gfzN9UKSIRdvpT98sL+anHpOSUmhFhlFcLs+Tkid2uCouewnNiIl
5754JIgrFb6un8tqN4UJCFAoVTQ1QQDxk682tIA/7WUeSx2xjlz9/kd+sowSBNa/K+U+5+BnYuV7
5V/oNdORUuuL9TNB+99NvLNXVGSrcMp/E87Knh58y/HFitSyiejSlLLNAQrwjmtICHOo7pml5LFD
DwzM1jjboEmM+uz2F4Xq7/3/uF4MTP16dQRf+mWKqq83yhnt9PCvn38ATA5RypJanj7YGsaRpq9x
z64DdG9tJtJYgUviF3x0D+Pbz2vUDSBgQC7NiL29X93/qKt72tDx0MM7pz6oJtO/YtBhCeZKa95M
JrjpYEiCL3on3OcL0dbbAafKEZZKU8nwj68WO21o5p6NmNcaYVKg0U/DdA0bp1iJQkqcKJcPCgeY
ffB6OT8VfVNZAPmHQK0HQdawBBxpOz/ft7tcODpeIbiOwqoYkwVQtRS1gl6TVRBzqlDNOgka8RPp
MPOSOmKUVZKLBPi6mpfXC6QAm4i+fpyOiNnB75zvwUguxeom7ciZIc4JUk+cvoJ13zlJmz0/mg4M
a0NCbNKWDSk1wxidy0vMm6KHSa0S1jM+gpgfufGceOPtSZmo/ihDBoRIbBTovPaUEevc5KMGQV+P
3hUvW8v0tajG1NwgMG3LLf5qVTTwucKJ19QVcA7P5O/XmjfSxi9Ue5K20WhD9O28IA/UZ3sbCys3
a1fKHdgJTAuDdc6ggabhh76MMhIxLUzcH4YeL4EPP0dM+uh+mX0EcBCa2l8S5B9e1a1NTsvGh/QY
YRoQkcW7AZ5jcKvo7ToF904+CvHxyxKh6/WiCHAfg2hJT1xcpl3Sf0HYmuLvaFm7AArt3qdHBYAW
Snq1KvJPutfzK3+SD3/fUl0CGsH594bU/zwKaI64+tDytIdaZEKNbYkpz17mJ+FE5TXi0qA/cCzI
zrRv7VX4nodGQrbNIKiPere1T2XgVdpeoDZ4b/NfcMxBJqjR2LogkaOkIzcxuv4rXzCTfz78rNlH
GIIGDzD4/IIw6dHWIkamyBhD3YYuiMvVdFxPK4rZjE9G06PEAr2+dSMHeNItlYCDvBU8KVCF6jaC
BuqhMDKKmwATYesETfrO6olKRqFQEbxLJGFOvcZfJh7holYEKWNAHrrggNMXpOa+7qFHC5WNh6vv
2IZyVXd/qwtpa8fTLnuvFjyVYpc6L7VMCq6elP7G1EReT4nBxYIzyq7CCF7cV8ALedCcGTPz9EbW
PTlMrxFihz7vd+2HVt5IIWhyDhD3fD6+hL/olso9sLFBewoWBIFxVFwbL62kOcWBRt1TaET3gDQW
v4PwdYtBeUmgDbuqNDjHOYot2OjFU1Xb+xdhKeE2hDlDUspyqm2WUZ/n/qrJNwAQHlkUQX+U23wy
HhPwsqS4cL35wxhFZ7o7zOprNRs2ONWDiwiFRSiYdLugoRdgehbTWQw0G3XdO/IkzIdZQRqTZ4oi
I+HqF/ou7jDYw+5wWwOZN1vQvdb0CGCgltD7gJlmAW0egIcb/K9Sg0r9syiBKj3Gj6ffvLwW8MP/
nP9tTX/1kCVIvAqIjDg+IwEc+RMV1pQqHVSpB+g/aOcnKHFY5lbSOJ0GoqZKnxFugbpjMgNmZtG2
PEjec4xL7gRx6LAtFVlOnRLOzdHuQtlSrBJrewaLwF7MVCt3aolKnwJSbkr+Ig38mm25AxvLtrpG
JeLo9a+DfcSraea53FBYPB3SbFUeRSMQs8NTXtJsFhx9UnoaQBDmvIOWVzRKss7dBHCTDDyKds4a
SIWjyKHtvAl5P+WGs1m+K7nZA1tz2CDLaH6bd7Q6YoZ95RrnhsuluHaurbYgQNaIVnYPMxNL7SW2
3IMibuk4SApOhEh/O/v6hRmwFFpE/zuc2l/3tX+Gnu2C1o9mYd+LOzmUSdRr07iIo61IacicroBd
OOUYGsCh08/m2hOiEllxjylRWoU4xwD4uF/7dYQTJp6m2tE2fKwN2zgEjwBiS3pOtfzA/UFxlvEP
KTNqvO/UIVHwlKFK0yvRMTMSM/sVusaZ6hKNnSPrTtI07eKAf4Aouyq0oFKAb8wrEuGS8ZK4+2+S
w367tERpVYH38XJcmAHxVgZmvYhuG7CAopT6qj2CsC8xZwIid9gHhdyFZca0e5gQkz8oDJSSQ+Y8
EG5BA3MgCB315rFD91eYpbA44Zp3MlskX5xV0l3KTum2Ta7YzwMcIciTk2HuHtQiMa5CrM/IrmLv
4UYBLxs583BPhLwUk7zD9DtAqV+QQqrupnC4nSRUqx8mGQ/pc1uqqLhbi1FfFGN6FoLwIWpUKmIh
c80nW7OaZxXpiwMc2v3iuSleaFPNe7e28qNtL2ZtGh5hrsvUz0MR2MyeS4Nu1MAzROpMIOHdAFy/
a+yZF7vMD1tFfcwBgHAWEq+6anRQjyIOCch/H4zbXydHmlTFo9BSbEp8WLhxcC8XYO5H15T/L+SK
DgARZF4deZi7xr01HS6Zqw22Qm6YlFlAmwGr1SeoHklgNB8af4ku+N3+2d7zKiBbvujp2xD1wUD+
tAlwuBgL/9t5SODxUOLVn8DKa6TdD0KDiBnXyzBar8Z6nod5/rnyVQIZ5fhaJLo94ZW5pRl1BUUq
jUs3YvMfeMt03Pwam0bOKKFIy92P+CntvYcz0RNNS18bh/rDRHddFhy4wpLXIhaIIggNiS/Q3AZZ
9/eXfElclYvj3HVUaYmFzjfywko706BdHhiJDFZ9A0T06/Vsc+0+aENad1mnV7rr7YASYbRYKteT
/9WJ2r1pK9ms7zuTOtKDKpi+I/2N1lWAaoRKQzppkTRdJLXtqkK0cp+OzAcvQHwkIEYPA1QnCnvn
lie7Y1//BnL2PpX3NUqOmGvoDw1g4p72gFioHTbF8lmV/oHT3EmmYwKfZMa2u45GG9PMRxMIXYL5
/k3SDKzjn/EhU/ClTTgFYIzLKIPtcVKk4ocENuEchZKeHHghtiVhx6/T3UlpsbxQHGd09YINcDIK
syiJjW0yOPY2GlFYoWYraV6N349r62enoe8RPQWj5APicoGq5Bg6XVilId7HEz7wJUCCIn8+BQmE
ubBYaHp+3MpO4BPzf99Mbjqz298v1/abv0bS1qL/195nAuLpQoQgv6bAtA+rdklt5GjYoYkAIaeZ
HCR0Dl6VEOBewFoQ67J9LNgvZM24XChm7ggFbkLKvILRvUeQInq71fZlyCxjGpSNs4zQ+AZ7il4g
PxCMAT4vNU+vrSlvbCNnyrs9D/mEwAzCiKAKDziofEcSPfVilY8sUKGAFFwPMdt+0kAPu8OHK5GM
qCzf0ABc8cBCSJgAq82uIzyZ18rxEW177zTApjkEnMypQZdB5IYqlI4qQlQe4Lhpi5XaYtWPmtbl
kcBjuYrvw4pev9Ox5UQOHR63yquQYQBSEGFOuHJ6jMZoglVJe0gWlQfDm7+iWYQTzYbvn8ZFCVo5
Mm5X5xPiQ7ree07m2ZnLFmcYIYqlH/4ITGsHCoI5zdBn2+pYGxSYMMyX16t+nM+XKc6xRXhTovDh
Va99pAqRKa+awwUP4oJrx7I4qa5Qg/vav+wIQt3HulByWDNKrBhqRtHruOIoxFyXoz8LrNExxV4f
sb0JkMynM29az+CcdUr/iognf5+DJudszptBZTIzdt9ASP0jkdOdSSIdkVzjwzXVVUTEKBG5nonp
ZS7O90vgSqYmJ2rIQ+AOSL5s/2TdqWL30gQRdN3uEqG5W7udDoJmvXI/XlvBbtJACdxJmj5pg2Vd
/7pQe4v0w6YNoUD6ykSUFUN7SBSdh9YlFpbGuul/sV1H66Qqc688mp0Mo7jmPlGuxyn2IMJyNPkp
upRjeM8kEVt+VZlkoZFjcX9N2tfJIStGHvFuwxVkE37uBKSZi3zECZQAMbEnlRJEpO2yw9LIGtdF
x5LCQ1PE4bvUAqWrLMblzA1qbWdbMhpU86miWogBcRNAR0G21WuPIEAG5F3WMc6yq7gixww/YHws
1qYQQdeSvOAOm73Pn4wFmJCLE0K5izjhL/B2CWMF+HxFZ1MKCNdcpr9QNCUgqY8fI4Cqote9o9aC
kCihA1KPi7UGxHfaPZ3VjQ7QdmuSo5XqN6r9gKSG8pFzB2eqroqXR2DqiEk7JKBPX2w6PyYnKLVx
sqHNoBN+Kprwz8p+dORfDdGYGrBiDGQCsGfV9duz6DSdNBPLesGldNtiIw2xd3YzyADnN/LRSYBK
ti1CtZR2cw3gqQJSCqcKrglSV1Mb1YNBodysL8oRSfcquuMcjScp6TwHOcM6LXB4UdsrAJ8pFhr1
9QHpJtXjiJmydGI1NOTS+CdbxLYreg7QG9zpBcz/SkQa9woPMWTsePgSfPVws/7uqMqVyjUYtyj+
6j0Ud2QccQ1IS5YGMfY9wYvDyy5eZfoo0BC3hRBiVHrqkQkkDHKegYK7ds7YvBjYJY+zX0hb9GWn
JxFY6clnOuj+ybpg4nMdFVXg/fSpoecQ39pAUMJrX4SPKI9XE8CpYVyY4C+ysCv+MFPmoRnQUbms
tViWaNhz9vXcdCsS+I8z2hFgauxYu9+N2UbKrMldEMIgpG3bMwGifh98ei/HPkTiLG1xSpKwABZH
5/6Rha/0WuyquIX4HViTx/dJlFmXOunTF5IVdpGntJ/pqhKKerN5vcsUyzFjtXFRVZx+adxuUxZk
J7dX4LQG5cpJF2+2594/Uwiw/CCaq7w61Jsxyan9rvavpN/M+L1s2kgk1GKdHP0fvm09I+ndPhHg
XrD1wx0VmWC5+37imJ3z7CScX0yghnpXa2YOYBlF9gxg1+zBSAnoGktStqvGEDka3mizY2lRiDAv
a7NL+WA29EpBUYgbL4AyHraUF14DSPD1PclGzGx2AR8UGxc/pnFJCHImrAm0Umqo/lTqt8T21aPQ
0P6yRs09ltDEVQ0HKHFRBJxc0GtrbH0Kac+B2xqfyL2/V29eYtI6ypM+Sm8O0Iy5OdUpTj6KXovG
g3YBuo70/2UV2c7Ta2bQsiqlvTtFPL/OVH/oUmOo4OZAmlBT7cW+gcisa64BUT3VNk2Fwv3wY+tV
20WNlLSEq2EYvDCqcUdsaz4EA33kkHTL33utoYKkvyCroCG39lvSV52vU8O8B3XKUd/VewKYpN4e
8YR1v4OTYXvugNC9GWacovp4SLlh4v8BfRNcoic79o7TktSSiNw0R5BKT3L5VH0ac07UBmcLMdgp
5J4tLhR8q7GzMzkNYrbgvoX+8GDoya8TuJ39uycF0Q8xnMmhVdPtKaR49qGSiGuVXgKP5xi4A6ei
/CjTz8WKJ+RjnFrVyKfClny4wO3nCwh4uqctUORn/SVXiY9UCP06CEawi+EcHLSbXbu4rStHoaZG
WWcIlbXP9o+NjnH362tYwl+Y5iZDQqaV/ZREAHEdUImWRnVF9+HeOnDS0rEuBtpQ/oKwEwQ/PkaB
wZE0Xm0LK2k5mccWUmCBwvXJ7tmMbBjYX3ynxuGMbKGohFS/0x9AvB39rC9EkMVWnkk2RvSlTiss
xJ5C0gaCStn774UD/H/iBdzSLSWk653aYL2h13asrXs34bKe2vdz6souD5kCbUmTmYq+WwI4amxP
CBmr3WF+NlhFHqfO0oEJdMcXMcNO3DzfaBL0X0ObdoPT9F+DH7HZei+ukCB/qkQspUSThZtL69d0
xfENRvRqtJ0H8PdwFNzyXHdPkBr+I8hksROzwethh8Gt9MBHAVahpDmhhrN1W9mVccI3uDFkC5z7
fJ3Hkf+rj51+8urrs4KK1gLLTsT4B/1fZg2VsS7eyyS6JqvejLFulukICugPEWbvq/ZJtAhmHA7x
VlkJsj4q3lIVMkus5sPVLZ/nBNuELVV4ToWZRHa+otuVkdVBfk8whvUoOkgtEeLzjXcFByk1k0gh
VeCNcobIqf9koOFbBy5DRW8mqZk8+JJq70kMwp81jvFPWfB5N+GAsYtWhl/izJr12cPyum5TV6Lo
qKolBmn5GEliG2tEi2bESZC/mS+pWQqXBgJHlFd9FIfqX8zWv+4uxX+yRC4IGzmZDA6qwFG0ew1f
h+0zQCJkhPZZ7WCrfbRR5ZuhBPdzFW1DPVOFFSUp6Kvslw03iAZD3yfp5sguyIqnLygWg+XOfHT9
ueXCJdpWlzro2CBc4uAfwbAvtl3eqvBOsBUvAs2RBtfCttAQJqPYjHnjWLkj/L4IuJNLTxfMZM+N
QLM6hvT3uRLPhggOnpJW+Dp3ki4F8jWZaDFxZBPyA7b2cEpHmA5wQhk+pu0sJREv/jcPH9jB3JDf
M2OhMnUiiF0feO7HGTMOWcc6kpZNXUoeVz6M5Pe6RJf7cXoRppQfg2FAiNCQHho7sd3J+61sRQi+
eO889chcjk59cQzfyyu7w0Tqlinl5R+4n+4vQkqGvY8Y/icfoZlB0lM56Oi8NnJUHdQT3s9eaKjP
CtZSzSP5nZPmQKqSRwr6N3fqhskefhGDVLq2HOSfRJ2brzyNemK61hf57c9+zahyI9CAFWXpfSzr
Op3su+d9krENcVZa7rkrXIUn6XFVAPJ7cpYQuNAAsHXJ9b+wB5/8Dn57guDewVqYx9Fl6d/dzW+l
152ecH68FdYtNty+KlDbeRI7JdUb1ACWnjYQVO3jQfJRL+4aPm1kHo3VgQmSaozqaVaB45g0v6hn
KAJYmxHJz4K5F62P65YI7x9SGl2RyCRy5NYt+wI59XqfJQR1zTEcE3QjYqwiafEiK/OOpA/yY8d1
/t+jI1NENPZ8YTHInRAsEhgQBJ8WX+JU0yUgBWy/dorha4lE3IFUXQd+n13kphpPI04EcnRWBi/g
W+Y1J4TRpfnZG51g2CpAQyjWtGG15N/KUcbp96f/es0XTA6wCPsMvQHPnrHD+Aev3xdIWuEJJN5N
+Bno9Fl0aPDjyqIAhK2No7cg/zXx8NCTCAwIPpuUnainAoF/d+aKyD+g6zQjxqZP8GSEqrKsvUHR
QQJxsCCFZAgQHoE7HBahPa0FJZ9YApp0R5ohOgLCyEiOJQQwMCAU2Q9C85eYB9De1aePn0fdtM7F
Ktm4J0wQqDKxfBDtOm43YgS6fYEoVgTH4GpDXjdi1of9DHrmwg8WWmHdj1Xaz+8MdqF5Isy3krrj
h9phv0IdhPE1j0x4q7JGIBGj9bzeMvvurGqpD8dA0amPv+aJOd1t1GSE3ORiVt1fqmdvb3pAAG9o
b6lxHPMiRIeIX5YDDoXBcc3OQ+4HV6A6Ct1UVK3CB61/yzg/I+OwWBC/XgAP6nNvOIIA2KrZv6fq
gYIcI79LPsTh2+YhCnsZtKXhX+/tBKZpv1wEgv9OJATlsEMGhuxKYZKX0rgSfYcoo29skjfz8LzQ
VNYeqPT2A206VRxzA24HH/NRt7k9PkK7Kz0N8JOmUTcaMxiP4q2H4WSIfEk76+nKnF9XfnrXs95h
uLnTZQM3li54XzGx47bO8ZcE76MZOlUBX5H/iktv/I+6hRXY802BmGpGW1mgZtp5Y5YatCu5LH7o
2rZjmxI1DmL8uzX31iEGcULeFlZe/jh8491kAo+wf4uwq1ELmyM2P+me062NBA54/oiGQa0Ig61G
l03hFHN77F2xBMiaUjdL6lL5Z3fl8Uwbz6K7WY2MzO0YvASBen6Mi3aoYPDMDaNZC1/VFWtnZ0/B
rs9cVtuQjrryFv2n15Sc/7VuEkp28UaaWz7WXm/4Rt7z4ymRYIXknmd/yDJGOUDDeRqbRYNAOg7U
CFfaXkArsLF5KvUsfxI8IF5YxYBMeVCGzrPPg+JHnDkoX7Hyp4rK+ecH9QxTy4iERm/bkZGbKW5f
ChMLLMr06zE/pTZfXfzgx1PhKkZlOdN8HUH6aSVbL4P1wJb/c6SkSJxCrvX5Nyowga6zLGvGqGWu
7JcTja0yoCZjxcPD14npnUrNcEdgI9HVJwCERepPIzNaBDm/5kWTqG6rX80wRx6O4EKpH5pUt1I+
0lhWczRdbKKv5IJE8xQ6GfckKY+JftUrgBk/hHjwNLVFJemVlnUd+eFPeA/Qdk4ND6REQlFasf0h
1G8xyJkDRd6/DkY8wwfV7HXQElgGmPQ/toV8GcZGvbLAAgMVz3jBoITYRNhrz/JjOlgEZV5cWr0R
rMno1rNzQDUBzDb74DFjWBASI5M1Sc6QjH76TIAbzoO3q0VDSCbqluKcN83aXHXIExlWgH+MvqXF
BBqTmMW4Y+mRrFpHMhme0ZNzQEslcIH11nLOnij+CQdns+oSuHHLjgvfpDFFHRMSXjoG5zQ6qKHD
Pq6H5VxTq+86xpDEkAMgKCXXNEbgS3cWhI9HfmuShyNrYwbqEhcKp0JhlX39Hl8rMHekrZZRerfT
CQUVk8Zh/00LLRlRyIhdL4QBbiZMx3vpM0i9as/odM51VB9AeHyp1+4VyLIWt3m/QYz4upAidrgD
CiYSN31rS56vI7Sl+o3GPXr+bxilFTFLAhNk+noJmudQV22XDXeSvvLU6ucg4pt0dKqq6ln82Bit
h7tJ7SojIe1QgjX+PUJGhVegHFhyDq3pMf0fG/nuF7+AtEpxdL1TLFMCmRPdcD6MHKAzXrrX4sLb
bNlx8j1SO2s1/ZmOrJMqbMJBxRlOdpX4qASsjKp0MEpP3oLwqbW7Piokg5rpNGRSPu1iv+W7RuQf
0LXRoCI4Dm+jEmCaei+S5An+pR6pDtfTuk/U9n55reT0WJQvTwhHNfyNZOmONsWTxahjYikfNgJI
seDD6PLhtY/6fVVEuT1NTKtGWFrNos4tAZoqSx+HbhpI3ZBuH+W9u49wAklSNbchrUY0bE35p4si
h3PCDviPBvyXnaQvKxy+jMbfd9D3fkJ7Xwx1wMaiL04x1fh4KME2wlLZM1nd94WOcBZLE2c458VQ
unC0WDi1jTpxhcfNvsrjiDMnksSmUWyNpjxuhEBSaOCikYZ18kLe59FC8T/5BXb3shvokofdgWzq
BB2ha2UJyPoHOZCMAzh1y8UKdqjOrji5NFxtJCzUTCR+IJK9XbEJ38ebYkzLZkPnrt34MAy/U2GY
iVqhXXYUl4evoInI4Ix8TxVidAjyg5xQMF1bvFPtWqP1YvDdt5sru1pASZUMXQJg7U1h9qcpxDTJ
eawy6SOXyqv++s4TU+DDwpBIDfWmXAaeUpOQaYsBJROq0HQl34dp4uHMWCOjqbKFOK1yMi99NRIL
RpeEY9jWBzJWxcmPA3UtVhLQ+DaA381LTBuirjGGKIg8/skI9gr1QP0w48XD143LJaVe90wLFsF4
tOqzxtyVaH+vDwvBJRDBYYMYkFXbcqboUMh7dopTwLreb9US8FjnF4VcHeKocP9C236/AsRAT3b5
nPrYIFzGQLG3i48RF4QOyxTLrmKZrfmVCc5Hy4584hKiFE1ZpTMP0jTxNQc6S6nezOGJYe/f5u1W
dOnbTNO2vHiW2Joe8koJip4PZNo+8mduQp5B+HJXT4vKvNLjvTRhZML4Lhn3CZBvhEOLIdRj+EvL
YyCUlesoKpqwERTxK0rZvY2tvMcv2RF95sHGCXoJRHRtlULrb6+Dlso7nPEvPEkOEFWwGyQfB17m
vhJz+tNWWFevrRk20CZk0O2K1JVcgNyFttzss45jq6p8NmzRjFQ23XTIul7iothqYHrG/sXzY7q0
8QX1f0bS6cYsq1zhJDY1QtKhqFv4EfYdFqrwug5En8zPdfV5Ez+M5nfSz4EBDUkFk4KaXCL/0AL8
Yj4aiu6/iHaduygTcWAVapNcruAQyXXGojosNXbbNBCZyRNgare6ilaTy/joHM9+UlLAenVNMxAe
A2T8QzUQilbRxXE9mN2gS7AwdDWAXCB1m6rs1GfrkoVYOOt1hoBPv+r40ifCECmATgxJgVSZ3Ej4
N8Ud0edeZO+lalobbAzPOlArPaHRk4UmLRTRyXeeMF7N4xKGOqX0XaMFfGT7TQl4nEagUIiWAoKV
b0Lx9MyVhYplaMWsIxd3RM199536bhaTlRhuUHhSY5f9dr9YGD3fNL1zfd7MKJXa+dleJkeNDHKm
j2JzZJqicwdIDvJH5CRQWLjp7unsfKO40mrf1efWj2sj4d2DJPjbpKPdkFn9aLyW4FNVw3XKgirZ
gsLRS/l2FMGP9gSUftUZR1I7BtIj2fHbP9tgzRD8uuPTLNb6hIUMZvgfeWwPlREZFQAkRYVIfK49
JeAhnytSH+Y3RwSMwiBbXUStptHF6iSOpG4t4SgoU5JYRFMEAbIGObOHsfbEaIXjiIusncsT8YMI
gEOHntODlYvyBLp393Rq31Z/P96QgRWaG3wPJU57pAmgGNuV9co3gix71i3JIJGcWtc7wCr7DbAK
zycWL7BE2ZG2rgiLzbhfqik0zEy+kvMnhNUNHmroMxlDM0vI12UdPSNiuCG8XpBQFOobza1fuzMu
KDmRvKU8JnLYNK+gW2rCCv/dOyOhWO8bIMtW97EkaA0vm5caln3+CbhBfzqaJ56CZG53xTZr8Aob
v0whChbT6TA1N7AUeT276YHQtzDHHlzmzwAnXZtQfCr7VVo8LHwt0wLptSYgbqt3VjiT2rosvXOk
eQRfcfXIWCmbWEy6xdKGfBws1oho1BsaNHjbw1DS39gGZMoYoL3zMGvCHXHiq/NblIQobduUahyx
3SiGkSJtj8bMUJJOkYqr1nnrDelzju87DVIDKzSsaEyF3ckdSIEzUBMLy+wBFeQFCnMpNVNtE/qf
dQGpqoubbdRTjObYPVvhurztwTGBpZIRlX0Ghl6p6LwEUe/ZW4AGr2DLb3i3mXQZLAB5Eg2jGRrS
856Mbb1EjT+3g498u0nzD5vr7xcj+gxKXqqlJa57N//IF+KjmajRzhA/jbGPTvMQ3tlnJSYt7+ln
1QsF9VBFHTzNaee4bVGgIXwSkEomAZ8lxevojYniST8EgpPtRcFhPgZSLI0iQZhqQYcV7qoOhQ3q
iIBHo0fWKal1wjdEtEL1XJWGGoBsLYIJke32+Rke2oXa/R8tMzzUefO/r0RjoGMQKEKFko8cG44+
IEXd5AfCeB3i8LspsVXPcL3YmTQPZKzHWHrc22+UFm/IcHt52dyGmKRAV1rKoY9qNMF+vBUBXq7R
SrWFo4L+GjvkjqLikqlChHs/O8K2srqm7m4dcuEg0yhZQ7XJQ74HuAGHZQWbbhuQMOofo16ejXRM
h+7ShJpl2rFIpzIOmlYG3LJ4tx61ChH492/8WcGKKZ46DYAkRgAREL+GQdNNHp1QO0KKdMn4qbwR
tOmboeb6PtRfz9cAjuSgqXdGNHd0iah96VWIcJV9vlFqj3suRrtLixXMZFKjYQTsY4Xxl7cVv8pA
+AjdT+YMAxsw4Qw3C/kYnaogHAPNOkk6TappLCtX89SM6Lw52xvKfi+pgy4GZwov1UGuES3I+eHv
8p8qvdEuWQxxNQyF89SVoiXwQ74MR+PkYjmf6II8bIN5yGRxdwOOGq0eE3LRDkK2Zd0/+J4tfIR7
vahiayq44/EdUveOtzu/oI97CDO3Dsx0lc3ntYWJCZMDoB2ELAoEorNw+kTKEXJVbtJeRH89nu4S
sdbj2ucrrszsJ6ZFKlF0KWed3SBO58lhtmPqOZ1WWuuyCr+eN4Wi/m1gdeJYDK/CmF+Zn9kg0+UG
5MkCCT5sEhA7kc5bQ5g1bCsCYgXsFIQlerLAsxosu2eM7axSvAkl56ML7PSu6N57EqGsYzWMRRQU
hCjzl9Lv9IdxJxG3aSV5OYcJB+6VaEPLWtjmPY49Nl4J9VBeKk8AdjJjEvHMoZfsiWbUVSlo6OMS
kuGmS8EgDH4Zs25uuceKnSfqnh052cIEYKxQq/ub7UJoetS65f6IZPLCzL1xIOSAZZvscxFxi9PF
aOLoE7Q7D2hRK6/irBLnLeOjRlahgVzCFKQML+xTjkv+KJYOcFSHRFF91YskQhmilwuT/fRVk9Hw
AY9EA444503SawYqIHno2tPNwv9ZO56rXrBtiZ6vRUqMRBLVtjGTsM6y3UG4KK+Z/dQDiBRXhVKK
nkF+8I00hVK/6cVs3cS2NfLYh3r9MNA4uoMrtRZwjB4BYTSN/J1ONgxqeKWF5ykHUg1qS8Z5CmyD
3zOxp4I3J+6eZLgwfOCSHMjIpr3aSR5485Qsu8ofrUaaiRk9j8PveqovhbqBwbgQGqTzBjuEppLC
HXofT2hL9WYTtpW3DHsm4vEvz8+UJycSwXpBayA0qCA5phdWXENMgmFDkYf6bc4+l5AkktGvIA2V
rkT4y4A2a2XzBPehyv94ygVveRcisK6WqAOTZAIhLr4X/Borpf6IOFeWIDnt6b89UgN6X1GVGPbd
DfLd0SCCe1sa7XdCUbURFuSbfGjfNhVqK3V29W6sQdNdInloNtW3EaGvWPA3IlaK21+9//d27T+i
7B1S7yeIB0DmtvfY1FWG6M4D6v6yTCom8+F3F75rPwcJ+bqkZM8jrcPhc7Es6fw1gc4E8WI1Fx+2
8kMr75ODSDrwhzRk0CZ+D8pqyMTlG4qRFavnwpTc3xXx1ivVRijF/EKkEzl4gCDfNZ8foP6ALAzi
+5rLyLmOOd0gtuQXpaH4wI/l5CluTEIgPSAkSYvyawWc/4hf60qxzCwWlqZafWmvTxpwb6hDitVn
zZ/JJ75La3timNsKP7ElcT1RXU1Z2/jX4awaREkOW7a8D7Z0iB8GLxzHjhb9hKt8L8OkDeZ0FB/B
kTvLo4W1BnyRgFl0bPoNqGT3yYtpTo8y/M/5/KMUiSc34yXVw5VmQ2MHIgxQRHtBYaSsIIYPMDAF
XladUxMIBKCoIK/a3r7mU5Ns110f9ErVrBYFE0Lu2M2BgVHVRyCiWTsbx0MtSAY4vPtJOuFJZoAI
L0tY6Ibrzyr809WrbrHHMwnfsFDcLfSVC08JOSOB8KV5onX3LHNRj8i1AvJtuTY0vlI12Amo9AOV
5SHU+qsoJUMBKCtQDQ5SAjYIlp5xacwLu3zVzWIum1BYQPeGmbULWzSJtdMUu2r/mnmKz9AudXxI
cSZ5/KrBpcU96GbkSc22lWEfhIrDpzNGT+477RokWw/5BA4lq6R+52p3h6jWtX5LA43ACeZTvopy
BN/dQHCBlW8oNh2WrGvEkTelz6qZUkf3hZ6YIWyfs7+g1chE9nb1F1bnRcfa1q2r0t1Sq6TD8gDm
ilrH+iYbaM2Mtt6uvkRex1dXaW3W74vikSz0T+dpZouoXPPYR/v6DGz28fRkqitfMl8Pwy9yj3OS
hPO9b7DSxgpoEeSCTeETQdgvrrK/ozImt02YrMopMnppceC4+HlIYbJBqJvgSlx8duEycdk76tE/
cX3+yUUMrSJ0ZaELe46RwAfoW4q6igDfR2cJzLgUKJazfcv+rqfF+Q7oZdJL2ChqPO+AVCjK/smj
bUYWA2kfFnxaXs6s5o1X9HvrqblBzewXu4WksmLPwZ03Jwg/z7WPQgeolrQo7cU/tzOHgRLZ+L5z
wMU+h5CFRTl71lHQqYZ1cJmQ2OApmqFsyTJ55+8Zn+B+P21kC3UNACVYT+uRo0YwIuNn5FQgm5Za
E8HKGMwtfm7VtW9pdbsnBwHV8kJ8Fz06BTzfkaUeS3i6fKB43x0x4feDsjMoC+PoW8luvMpd9sPy
jF18abhAygTkeP653TZj6qkjeP49UAbNmurNAHEEdtPtRRHHXVlipKTs6o16O5XW3LJm1JrydihX
JZ5R0N8QfoejIxg+nq3n/mwhwX/zatCtON1W4T5DNcsOad2oMg4ffVQ11vTHPdsoFOs8ucfqfveI
Wci27BkDG+lxkTvp0fsA3n3aDDXP5n12pd9tFJbhD3tr9rS+xunqo2AJKDTLqPmjjUsO8KNWbNJM
yz43anAumfeD3/riRWa3HIX0L3FdI5df9IITtsRDZ4iW5b391zrQ1ycGQd1krBR4V6TEySH2Ta38
vIqaGzRKgC0BliJWCpImq0IwsH0EIc1hiePn8r9zPvuEbu2pyZw+sRIiyUHkLBr2TIf0X9tucLGD
jl1zvMCCdOrGk0XKcFarVFWhqhtvHYXZisZj4NS+M0z2WItn4HTuzo/jXdDKF9LChiWR0FnIVdmn
1do0yV9O5mcU2gEgJCK5I6bbmvWlA3c0gLZGTtlNRqrvsCpbp2V/2IX/je0YjdeoLRmyB3ETwGx0
2NdlYSw9wzBetsQmBUD4VzoJOvydJ7z9yQcWHKkiiSi0CyxvSqAMwMgAH+dzaReI7gYpaFsWOmQt
XWEFZbfEMENnZIGyuKXALJwXRth/CgEtdm3/4swHBc9NeVdoqfM9qIf0ndYiqzo7OMKD8PQQghSB
FgrGbOg4OQHpjSsl/rdEBusf+4S9jjp5s19aYSSxCeXB2BJMTOWjNE2+vftxflCkrsxmv7BL0M9W
lBv4R0L9YCYUsdUJYrHDQRxo7jAtwVbkxNjTu2SMzgRbECix1Sy3RvcWNkkESjxUunzpwHUs6dMl
xughTU8UFWeIj9OY/gc2QIWLFqHS/2HXEPV04YXxtIg/vLZzpZDWQQYqef2G412CnWjziKpl8gnW
w0rZDEs/+DixxwyA2I4oDVp+ThAuJqjBLkEzLkcrpApiPwSJtnhJ2y5UcjDqL0XjrKXfs5MJFPX7
C0zhE9E8FxK8YzSd7gGbMkTX6ZF01hWRMYyGKXWdGkvBQqvV7v0WB5gLnIlIkjj8Rz8Ti5l0Oo3x
IPFl55mJbSsMuqHZ877H9htr/H2m/WlWVknojg1S+xFTTs/wG0zM7+fL2CNxw01yntMYDwikrjox
QcU8ypRApYi84JkcFCzGn8CGtkt1bASCWLD07gp6V+YEkNPQNUOxtFKtJ+/S4kEDLjNcLcpWlQ04
9E3mc8uxQCIvNMpRteTJGgrY9sShX8pVD9VslbIDiiqGtE2HlRUcjTgCrcGhERLjkRyHodgJArJE
eeoiat1Zyow1z17yRCKW9DxN8AsH9CclB5BI99EsQMM6llIMPsIwxhWL5mZ+XGPB45RZD0+ymsi1
UtlT6lckoiFQRgDe3xUqqZpBgGpQeV5+K5KIRz3ksr+lMa4bP/xBiv8BpodXNYENzCJnMh8VQN3C
kSEudpIAXhDqz+vDCOBi+TuhqtaWDBtu91JITSpvDwRxVhCAyKXaUQmjUR4bSVAiELWU9idrNVR5
svLrVMrKpgxKA4mvCT4W1z7A2ff+tEDt+8mVBhrHHcWkK5cjWMwA9sH7WHxxSWBCEI3uhKDRZ2jX
gOpo6B0tlnSMD4z23Z4buQI49u3E4KYnuy7E5ubR09VNRMGSqUGu9ewSO9c2Gn3Ps/HeuUcnhqlG
pMdjVBjGgEMlCmrWX1OBg6WopEBQ9bkTa9EAMNvor7ZS9yzRLUXphHkJt5i8kw8sToIXA7DBrTgk
Jk5Qgfje1PJa7C9G56xjhh9m+SUXLni8afOYvLIm+zuRCp8ZlSfZRbvJJsuQ4XopqiLWwW0Kr86l
qSfEHx34jzQp4dhclQJTiel9RQ3NdVZk2821mAYNqIscHrqiKDk/v7um8jaFbc7roVCx8v6HchQv
ZLyvHhWTOir/LpQAyu7GORTbkHG396oeRvFePLql5h1fH6DA6v7fTn4w0p4O5+3bf9mZ+AOI/2fA
SfNJe5w6bLbNgA54RvkFE0Bqk7EByKhdYwh6mqUCFbnjCitTZ6CsLa4zhnCNsIqNp9oSBOGIhMPr
U3BfbOI0Mla3T1pC9D/8zsU++o8G8wCQWRQNt299IYHf3okhZY1ha7ptKrgpsHyoucis6KCuLwWj
Rp0mMcBrjJG0YqRaIJyk7Z1YoduKC6WnOAPEsbwOt7hQVAvywVZTibWrg3WW17N6i/vNDPQS22Dw
/9roEG1Zcn39wdsRqG//YwuiygwrBpG6xJgGIleiCxUBjwamXehFeU/6L+U1xq4cQJgmM6IC38VN
1wXphgBVwXykjlsU9P1Kx8dtCWpiLrnDC3J0JBU6jL6x/HtndOdUu1AFxJphuZSyUozP9lgX0Oru
uIB6o3q6hxu0vMGJL+n6i4+fYC5Ht159fI/IDFv9Dy8pAwcg1XLi3AResozqhnlILxZHVL0/FhMw
msvmJ9+Ujq5Mfb1Y9297bT4kDUQkaOV6ITgZWlHE2K10KqQ9HE8ZvFNcb/6UeRUOWGcLvU1lOp2N
b+RSYNTjWZzTNQtn5kqz8qGPcWRCTDnUW2VCX1EvCJurvMjWUsgbOpmIG+vuc5t+TnBJLOVKLhDR
HqwUCYSO2jVAq7Hw86+Kz2Yg/KhsEa51OwCBEZzH4qvVVTeyV+Z7tonJKGH+O5YVc44qpzZTW2uW
MSHliP3yDz04wK1rueIxkhoZpt6wivrvYLCRqcuMVXx5zhPTIw7IEuwNZcvoxXrKa/vpfxwRYHEJ
ScCAeReXISRIloG8Ic10ASmnw3ZcrLFAzexstf0xCNkgPTZpAduE4ZQFUAZaTKKwq34V0rnwKTui
xxbCHC/pBDGlqW0qmW0IEovGYedfuwclNQHFy/X3ZgUsnvowiOEdzEpJskZWcfoqiaXRbBoNJJ17
WNkL/zhavJZn3spzuhUyoteKCLS520bJn4NQrUm1iq36lQNVdUe1IFJuLpl/Gsy/7C5EmXiL/Rqo
YW5v59qrDBihLBz953zzz+zh4IH/jU6lznYYIys+julTyfIXtmcw6+eDCRUzXK38XHgmVGY6Ee0h
6fQlHoR/3RYOHoYV1j1IRFksydqSSfjyB1nN8XuB7bexRBqgZgB5wIBUMFUyWswNvl8TIfna+TSl
OqkqveK/8tNL3Yqg3RoPM/fc+dOhsOudoonptFcFu0YOinMADdLkYClNNLVIhGzDx1qTRm+2STwL
GPo2seKL+38Jgm2vuEKTRwDv4mKcRngax8abNB1EPt/7KORSsgbEhPLHoEfFrwpTBglTorGHkkYr
6EWKEFDGBX2gvdSJTQXvYgBqOH329iRR0Pe4dIOhSmrC7MNAI5oZbNyjJapk+4Tj0sOa4YuZ2b6n
MeDJQ/CSSuwDlFcxxVeRowH8wMywLNOmgIVCyxFZ1ZnqI7ru6dDun4GmR9IuNZtDyMeCxnQLpbla
3A93W0pnaAuiqDEa14d98D2NrO3NmGnsIMDP75Eff1heg6XJR8v+YYT29exH8NkUHVBpPyo0Yv0P
Xg+cBUVO6YBqJOJfgy8K2ikETPvfEHR616r04puKKscxU/wwrPxehZ/ifRZtJW0okEhdMlo5SAvL
NSJQ0UY6hZWtj6KRdPXVf+tC3z8RRj/wJsWuS4SzGMffpQASqfiXvs+Yb+szISbHqOsUS8mlqkO1
spWS6QYxR05enRWCbTuKBPOtisRao2Hzvm70Y2ORYZgddaf1rjFE98idC6kONvJrvNA2+oSYyPPS
+kHgomQji+ODXru/qnFI1bf1PW7hA/E7NcdsB0L8H7f07/TaL7ZFuiNYeRqIgnSq/C6J941CqMhQ
BmHXmRs/pdxT96x2/TWhwGp/XPhBvPK4WvhM5wDbo/KjXx/E5ABCBe6aHmQ3r+C5OXvN6K95nJYr
GljCDkwrtGKrUvYXW9qumRYu9STiscr9ntHGlQ/ZneCI+Gmjoq57NUV3r20nO4azxlwAdUuSpgF3
NEJkrevkeHwjTDIeIRdDmZGoT6gObsT+ux3Yss23h2yqrqrnwmjIdtq867YjPkTH+pEUeWhnRQ80
ddO5pZVucIUVQt9R+nQDP6tmQ9IzR0CPBMwNvPEorQZRgPwBrVJhsC1hpNjy5NNWJ8rsGOinkYEi
hhKMX9Je7Ajg2LkpeTfePrAd43iMBgAWSkk6t+FBH9mqFjJrJ7oUHEAOTbl7GohYwV82/83Bywbm
vtiyBMPAkhLfN7XRBQaP048YsaYCVkF/kf+YAsU8h35+T9gzZLZlZ9zZ55ygfgHTZJjUyc8XYnt8
DTJbTD3FuWvrI87lA8Ipmyoio01piEWux5jI/mgkOYpC7911qUtdAzq/tWXIkt2y1MVA88C2LPDM
426hgoei2iZ4R8IJtKt+8lpqoZCsHfzAfpDAn8T9Jjv0iA1FmtP2IQZawKafv0tVE6Xyu00W4s43
1WoNrkRhjvBApOI/c24B5MCQRHkMULpl4mUY0iSttF/5cWVLtbSiKN0r512rPTHoMQ3YGwV3CFPz
9ZTn5udqpmi4x5CrldpvTboYOBLYLk9Rl6H/YbU0MZF1hZS2+WV/1S6XLyvmwfuF+IAdCuO8PQR/
pgO+EN0aK82OLisBw8JcinzJ4cWvBZW0kE053WpUey4JG5srhc01U9HPPyWdPzNh1v9Ciw2UZwRb
umUzi2BC7zyn4hi/BXhd8W6tOwzJDPGY5BinCl+HSSP6X+2XQ2vA47PQR00b1NMwBKUeNAv/U8FG
gt1S24U7G+/H+DcmzSuwT46zW3DIS4hFRTo85Q3f5iAOcou3ay5/zyj8UN+MPcRDLeHT3IQas9OF
RMFReeLe+QMVGK5DFXCdhwVm7h7PfY5CzTk/W7ucbGxBdUAyJ+2vcCqPlCz0OzQ4fubPG3Lzh+ih
lU2nUmHBGNa+yj2kkVMBb3ZqtPp7+7le/OfBEg3utQIDkBKcUcvZ0uxAQX7L1n/kC01sgbwrYvnu
bi3viVfMEt290XTm4ljH/1G+FQyaYVVvN/vMMqbKAbfN3xymXLywNTDhwIg0+7cMm5A+Lm7kB6Uf
DVE+JvZJ0RvJGKBgrldHFByEvwU9ngwqtZc+UPI+k7m5bNwbuG84KEn1TZh1JVVf5VQygoVsCmEh
Ao3qqNnHU/eGPYEI4wJmDVoPtqyf9ET17S9YIXscJKKV02jOwXMShcl2LA/PBLIraMVxpQFGA1NG
n8La4u8yxMcE1P6Y/Q6UdE3XTSs2fLCC0XYUFKEhTswa3pRXrlNlcZJ4rCOpQkgCN4TO1yo/k+rI
rYXsNXWTj375FhKMIsFRsXXlysNgW3voYZDRA663mhPBjDQvBDf+q7LxJxHPcX5843Q6zdDzIAQ0
jX7H6ZvASpUpHrJmTFQxGsu4R4BfV1RtTaImwujUqy1eunDl5g0qpPKNTVmgQQJ4shXAvtS+3J7K
zq4SOTadEoWyTf+TH9fxAvRFcsa0DGcx2QGBrO/zgDX32pYFbrXJfkqRlgOImkJkc0/ijvBip1Ue
b4PdrxgGZYRZL0GlUa70hUo2drbChlpG98G8m33ZmhDyBj/l+ua54+KidU+7hi4VZ2arIKRpZoJp
EEi+uMYO1lzFX11VHkmzhyX67aQwRGhDfthBenYGzslm8gJEt4AumWPNStBX6DaMQkrsXtYOVacK
9Myl90+8qK6JqAsBlsdvldm6vtFMZU/eYChhFr2n7RaSTeQix3pgZrNZepi8fEv4j/muTQKujI0f
0TVDX9lMBFhgTA4zMiKGpnemfvpjGLP2WMkpkxJSNs8+V8qsjhOuonlWemFkAAFzvnNRTRyu9LYT
IQM0eNy3ioY4ATlHrvjQHObeXWO3MOg2u8gVn6HrTwA/mQ6IyuBA83u9JH4lEyZ98c61GyomWncm
9Z9sqD/a43YpY2xWlj9VTVtIZ8hK3+B03i5NDozXQZabadml8FVS/WSp5nMzZCpsWXQM0rh8nLVc
FCiQich/U4uDxMsVHVhKkxUHfivqVQyPkQbAqAo4tlm/MDP/JpABVOZKFUPt1YYfb1vcJNBUN61d
8RVvIWY+6mBRwqU/ZNy6saL+OZuIXt+BIwnLxrxi15KE1SIArVagM30HWW9/iyVs28DIXel4+o1r
RxO/8DijZ7fyNYZkVa+AzYvECHPe4JgFZigAHNIQYncDGXN1WbBc0G6cBA0Q/ycBxNZQ8AdRHtit
m1Zsq6MUUw4e1TRCKpl+E+gAJ0M7ptTc1+6N+TU856CgID35A2IjVYdQsjWiQnhrXVafTMc7mmMV
32zSnA9MXhETFE4yv7zN63Vh3hhcciYiaLF1pC+3RUFx61bdYJoqevB8lRmJfWYf7AnDw+uBzISA
Yq+Fbb14VkcQV3Ll1IsqsoeCG+EbNLgYi0pxaK9AiSKokNrWvJlpZQyuud94eAP6WBd61RGEjv5y
T1uIvBWNJ4w9Wl+QeAEfQ+CXXc4ceUCYLStLpj6Dn9P/tYEpkSz/YEmZNGYSbXPoWnEyO0qImJfp
cIcX4lEbiiKw9fqJ4SZnY0ayAb2bQj0IIX7OsgeDuMn+JjiUnR6C7El9VJUuvH3ub3L4toawk7mn
vZJoa/f1N1QL1KhspILpksPME6WhR0LdbxTHHCuqowMxO2aCcArgUZyOHrSHJmUXkkZMLIXlJH6d
rq1Ys3WkVspDC0CvNIaQe3tbPdX9krN4DWcAFJZWgHFk7rRQoG2GGvhG/Y2UGTMdLNDNaktFnRP9
jpTyAr1MXHzLGfkshDIVhivlNJXvbl/76LnnMPU6JoJZhWzJfTDyPoWLPT9U5u6fEf8sdBzL+h0/
pdu05K9VlK8n84T9aBkx7p4EkM3Gq8OSFLk0Jrh7/riHPNqGslQDDY80hPlHapyrk1V+iWFZeHpO
KsSYaT/j0UKfGjYw9pNIlHFECM18f6/gDQNkN3jj9Akd2KrutMH3X2za/vHi8GZ3aRYUfVwXQfr6
Vph/PNjsX80oRSMRfMAqcyG8gZew3BbS68lvgmtlWSQ0+ik+dC1V7xJskFfkyLnx10fgLCGrpy8U
uEzRjqDrqbyudnDzwf2bo1EnCKoNnwWgeJQeypBY+UYJZa/14AichyE/6VpegQX+Gr7BvideDY1t
5G32to8K0RV0Vc171e3iszxgTFFDwheJ9Q3KLuXyqHz/aPWul+k8a0/P+pZdUc/vZFmJmE6ju76T
pDUzpu1FTOBx5h2Lfm3l/cZpyHLuA2nemXt5UcqU4e6MLP4xJIOF9XjpPN+ER42vnFHBMNvFUTJ+
H4JZgFKxeiqW1kS05aerhKPJeIuT1eHHl+FvRK//J/F/cWOYfazkGMtEZsYGF6IwxWoTYJHAVX2C
jrAlclbzzK5275FbQLjcyq3LGFC5pIGHIMuaK50irRmSkSQFhztPS4ziHYXSaQjoSy8s00kqjPZe
Zgd+qYP4jYblVYfTnSFJ2iP4Xk/2n/zRVh9PBGiuS/jgUV19FXtaPZMS6adSgunHNq4Sr5JFcan+
gTC+Ptbj1jlL4sWTkmZ2WpxRw4x6VQKGo4/0Vdm6PcdsAZrL6iNnD7jo7E6SPzTle/ZP93M//AdF
613j0WumDdGKEODKPXzdBBTUg420o5c4JNOAlC0HtytEOhsTrlJgRFlziOg0wcc2Ge+Zrj3XrT9n
xaZ23QmDj4mzdx3IWn9R+1uWAVxN79gDe3lkG/d31v/wTunWwSU8G01Q14QHzMDmaJoFKKa5iyCW
8ILModrWsM4QgIed2MAN+OC9xEkLqzjosvFp4HWxfAqDt2oi0st67qqrcjmqmmdxXskpt6pB/WJ3
fSBZ9Hu1inXhdIKUVz4vFLsORkADxX3j4AV/NfsbB+J3B3XSjeWkUHRXDvoNw50hEqqOBeOWZnj9
qnG+iuXb35+XHw8RxJy0l3KPXq/IqubdyP4dvuBW6S4PWcd1tHozwRC2JnwU5kdnBSnEyzaXmXfu
syz94h0AdKcg/9lSABnO+7AtlpN3oObazkR//NqFgbrnceXJFpmkXOL5e+ErSeELOcLOTf+k8/CZ
q9k70YEGKDKCw8gSjkJCUREKl3jQ7jQCgxN1FBJF9/2VCZj3H9GiRpIXwUrRZkWt9PHmPBboVkbX
rCE+RZdsSl6krenC/regh4/VLmvzvyM3hLeufvlbR6YbxLJAlBHLtlwdEF+ytYVvvupkV/95hPce
T4cZJM2kUcMOyVuRLlqysSSZ6CeF+4PROoiZMPcSN8NeHUdrWr2L7MnO2sx1dJ8S0qOcnn97uduG
4TfqwKbniFXa/Hqkh0HwMNtm3ySSr7rBnhu5bcj7P5czQ/gHuZLu/+4s1FFE+Ct6Rcof/fCbZ5Oc
R5izM6isJcIfAEIvojJwT675LZquMiwf7fbmGBCdVvkcMiXQNZ0cgcfnz+77zIwkYmTRRSfPrfzi
Ak5Y7KP5Svs8AQt5Rg4oN74XPbkrCAdi/mb9sFrHIe6eP1VqO2/m8YvaDvtS23d6baHf4V4FVPAb
iFQDuFm1/Yhpl40GXULhxQZUcTZR8sv1E6mHSm4bTx+J3Mh89wBIEGdH30feZ7KbLB9m4M5Kt//V
fbc9ngb8eRbR2C3YbU7+Y03MAZaMbOb8oyBmnnW7XaJ9I+C1dnhMyNM7CVaf5S1hLjt8AREkkRfD
JoOyshvJivFTjeVwEUoq+RGi5O1q0psgZn5Qr3Ei+wJSC4SRL+xvPi7tUB8EZTE96emYHsIfhxi1
ZtHAMyBidyYLppxkyVFi7y2JrGM3YNZptYHxbDhyovzVsRedGtJzlMYlq86d17G9ILVeCw/DJfAd
7WGNevit0hNlOYESkxdIi+jro+0e+eRqgChVp7HPG3KF3lcsNyk91XvWQO2sCZGWanr+611QzpJN
4McF0r8ijhsp53/QDzSckTUZJe65Bu7KXbtKm1Y3k2Ej6FOka27mFfyi6WbcUhh7ZGiYCIOwGDUT
J3GLO8Po4NlN1VP7BD2bduD3PYVCCFDWJIlID/VskiQ3naEy4mSwkPAjcs2iW4BCi2wJLwPw60qk
g1+pnOyrK40FAy0cMmTcEdo0KlElHqTbe95WudqBpbZVExsvj9/YWMe1sFrCQjE7g3d3aN+vrPpv
BCGIHTHurOWjGLL2uCehufXNT+mGqskoF+YfEiIm4cMe8C4YI6TI5wanTNjpOCCPDzQuBm0jbo3r
ZorWn5XOIw+UvlYd6QcHjPJ0SIPidITRKn+ndPUlHCsVt8BqUqkkRPgu1nBei4L8M9tJtm0mRyjd
VH4yonUj/Em+NmKl4FkGt9+LqEQF7Wn4fiWu/x1OPBwR9ikrLSQrXGkpffAL4xmyy5utoivAg9Oz
gCTOu5MdRc/bPmXxiFXEs4fPeyBh2qS5MhPenpa7umLbzsHqoqYWqSgKxQR1RMefwD2KcO/Yet+E
pvVH/dEJZQ9JO+S8oS8ZsAawUjTX5aQw1XQsUpv/HFCEzxWOauXnfJUI7IthLlsRhsF5ydXB3Els
fu2n7AaOuQm/7+dvzplgCwfEQYtOt5odcaWydoImDNHclDc90MK3fx48ZDImIuOmSMoJMwCdZ/lt
+KfEYJeNVQj+jpb6SE2PvbMcU91WebLraIGj03b+bbK+wyhnvJcPr+nYhj0a0HVza78UpMfdfA4J
qK+FTEbN+4NN6MG74X3fKr3PxEebGl2zNmPnUn94NONaunkxa9uGfunE+4X+Is19P9Gb9194UaEK
X98KXczzSkiGj2X4gBJX9cVV08knmWKXfytseiPCgcmWTp49wOPmXAeBlvuiNRKO60+bdbw3tMes
ziNy3Gb1z8FPhyQzq066WbdNnaXvI2m1TDxxaGKWU/3/nAfMakmXwCsjBOdPREUoOA6mxJ5PIV0c
wtrHK3erhVSF32a46zKnNVG9NNszyF+0g1nxCWygzOsliiLghLMzhxRLDXXcgDMNAXjfEzGLJL/X
lOvyIKndPlFkW2lCYck6yemWr2K9Fvbg28uwnDInlOOZtBCORMYVdIC28M93Cts72ioww8kGjNVV
RIVcFI2nr25lDuJZdfJUNfevQ0f5H8a3Lg3CUozVdB+3yry+6BcuaeZ2iPwDVk5ZDM+y9bnHzgmt
NS8keIVDc44NO7K/CnPL+feCDSEKEKJGbqLpljsFsYn6AC3nuNSrRmqlaeMj2NTlYEm1A7IaSvI0
jdLc2vg02/Ba6e9PLHtQHPPRx8seY76rBgA9oR1a23pKRfpDiqYKFYgQgBieS+IzvH35OpcNQ00H
0zlhH1ixBa1zba1VYtvJj1hRdjKhJiy31caZLwiSY1TLfVPrgPh5apa10/RyX/gKrM2ewpz5VwjY
7Rb8iVGYRbfnrywSeSQ3UA750D/UJ6M6h69dXKgTjwVhw6adJkn9g8ZOc3lNf2Dv7RVZWk9tPR7N
idIalwDLbVhKEMTqu3FGoxUOsVQaz8UVljiK9MqwB2cRwdDzyxcvfwFfk5+y3Ef795GOTk5cwcRE
zwg62KbSCQutnwZftXizBWcR+mKP9yJ4bebbwmRBeSW3g8MiOO24Ar1b7xpYpsNj+0HrfR0M/rP/
MBiAA5hzOcyb7mH5AFHSALxC1jCLT1wSPofM4N34TNMg9zHoqGp04y30AUtKy/Z54RQgqhN89yZP
/C/ZjceOEoO6/LGsRi1OpMxXJDojuxNCDyhjyei6dLK2qKNvSN3/1y1uzB4lo5f2R2VWm5q4v7zr
5X1S8j5WnIG77VoZPz+2TG4taggnX6pMPIh+lUCeZCOfmsHjBqERFzusddRTDZH8lsvwTZb9wa1o
Me9GgnRHr/FCFsfEMUBzAbXxTNYiFPxXAYHxCh1oFWoYlg9Xs8/L5j4F5xARW8VmjfqWfV6m8cdd
eE23asRiyA7fpzyCY4P4JkrBPJDzGIVeTp+QzqAK4opIGcQpVOYz/GjyE9+Ze0mrBCam3cGmwYWs
1eYDtN3C8bSFYsCh6ftYay49ItbBUhg/kElA+hbhf87hPIH8pcRMgaFP4ro3p2M01KR8Easi38wG
j0lDCY66/IOr4TMJunBnn2RWl3BKHyR/pjDW2I8+51CEAlSF84KOCwrFE/cj47VC9/VT4lvpzJA4
lqbZ8q9wktQS07tb+48I2u+a1dHbbKP9h8wFEATwCapTXl4jO6l0KFHx+yRri19N/BBVfUbvmW4r
TcId+27R17J3HcvGJ6HjXLi+eHTi7OdW37/REcmONujbtwlqFcNh5WmftvOeQUvxKBKEPWa1lf4S
xxEpzXreBcX8YMg9n6j9iHBsTc75MZdiujslugX3Au1GhUoZEAilmZjcSnyl5zGdtd6M7/Y1pPbk
EpEVWuvTxvGXu5l/OJ3IPiDniZPwXejHV2yo473WmFqdLdjI6U5XXr9uAiNzxUBrl0/Wd2Bs7nLs
PSqyextmXhl4UNtfQdkHDIdK/HzTe2ABkGOrCoe8H/k1pvlFqyVl8iTDX01KV2dtZmQVYQvphqyu
3n2nikIug2Pbq5K3iw/SK2KSnw4Onc1ITn7JBpeiJONlDxZhmzTAltZquEe/0oSlFp6oG2L2Rlqw
o8vb5+LmkDaWmUdl9JCrUCSnk5CobJbGM6HDt/HUJhVWqCM78p47XkjdyShPblI9Px/vtI30Jgcz
ctWJprLTjfGvvrac8VGl/R47G5VaiqTdqWFBRhplnX9XhOYqhBohZP72x1Lqv5HuQ2xwFDsGT9zU
ah3Rd8veZTHwigpM2hCh9ZBzbuxBntTMfn8/3F7nOT/RzVnLC876yj3+3hzdxf58AgIdZnxux+f+
f3DypJb/f1PaovyrCT3ZtHw1B2yZZifhmGgwW1H3bp3cHUm981AKDQVWPzsP8AfHr6URIjhtpoTm
p+c9AecJeANI1CNNptWhrn+UzTFusavCSa2vj1/sKvZVTjR9WmPneP7y/T0gd7Ra9kb46fLL736R
c1aU1/wlwpaNkTOIl37IUDREwJHGyRnCPNvomFiwIxNf9A7K+a3VwW8/LL1W3wxcUnOeubp87icV
txVt0XdNvUsxTrb7To0WY8rfgauEv/D7CptLve8i7cJ9sZCVyHmI+Zw/PRxPD0cw1moC1W2CQjVR
UI46S2QMDSdIDhQHChVXfyPdp9Nl36D1Q0ybEkwYwXVIya/MPLF2u7kxv/uFRd0/bR/YxRRPwKqB
1Or6MgqZqtE2U189wxrwLLtSSW4m3cqLEhU3L4eh5MkCagJe0kLWG7A1Fz/Sa9z37erniOFIu9Jo
3oJekQjU8bZoWVTPgCmczvsby5ckO2qsioNKyN+KdvMnXfzM32uRW6epJOapOe9GmB0vfASdptNA
9Ox6wL89ktHvA/m3G38h/xy54bwMzxy8eMQMZNF47/cHIIVDFvUYH/JIA2PA+SBkvhkls/pE08Pr
QTLrI1I+Aa3q0E+t+hGiiFclZFNzn7P/iMjiL+7x937qHelkeuUNpb9gDjASbUtVZg5vjZUZJWMo
tawATbFI5hWTeD0Pr6ImBODhn3a+HY2gID+K47dmDNEPO9pTo7sGB73/JKEizUKqWgcPqzPisuxo
Y7TUkzw3a89X2CiXJ19S/7n96SuRX6X4EnjA8FGh+7COnlxdLhksAHgCKf2TyuIGvE7TsPLe3tJl
3e7eMqLq226ULzJZEwS99um/z3e+0tUQEF1AkgfCy+aGpSdl+wIiDntJo0vDasAXTwC7aajlGp9u
8g3DnFcp2qb2S3NKhKuBa9oi5OR6kI0+wamVXVmj7DJ9hmSoVPG48Hf8GuGG7nNMdQ18hPJ55IeF
5MvqYLgMqYySXAj8j4lnLB0r6VJR7001YQMTRKllxHG0izgIYTWhYoM2S2dxkPewhr22QIw4nwM2
AKN1BxzE1vEelOscnbb+v99DWaO9nS7NhIgYjiTR3nS8uhRY50zXlu0V15EY4RZwl0F4RNT4t00M
dYt3An46fAo5mV/gTnYcdUFhx69SNEgY/7n/hlEYWC2B/uKWliumwnhWXP/wEGvGQBGNLzBa97/p
NcY8G9nzQmBHIJ9O4vAOwxhTnIR3Q2KQGav8jocgn/75/4FBCOEsBqzP9vKdO6XiZTbMwAeDX9Qm
VNoZCo0XJAhhmkhB77lTBvE5tHgW+JSN6CZ68aCybgsdpJRmYO1Mw0nGgGNepflqTW3Sr6KGj86x
prDYiRdwOO6mBz/4SEK2Sro36WSAttrFRylqFVbo6nmv6UMVGIET8UUSF+v8BN2T9KtBDAgjiGFR
RbGuwwShp5MQX2ZeLg0GdTLqas3hlEWSKZIV0o8lbRyWZCfQc8g0/x35LJRWtzZNXAqxBrd8FoeH
GjMCkS2g2rbW+GyK3qlzK0V/Cn4s+E6DeMvpeZnn9M/wRsJQtVUcOuL7p60GU9VRxpHIhhWNWIws
yvbLBWdE7+zajG+Tz1SwWTldFMwpfd12nji3bdlc1DAc3WbKF0cNSEDeV0r0+8SLLFMXZ4Cfpqrr
NmEIkZc9/CwEWoOiYnI3D+ExoeioF1ivYE9SU+ySAvXAmMg6DjmjcyPCdvO0zRYsyRoDj5de1U4x
/ce4FzVhODiHkhf9Pu6bJRFlgd45QrmNJJn/4b2kQJYCYuOm8ZDjYQrjHvx4RAOs1W3hO5NheRhF
5EiB3bKMOoyqePERN2z0wfKBSYOZqe0NFd0tq0vTG6zmzzNsUhh+6BqpeygdU3qqzFjU0p/17N0i
64xCiflhUwjfO911hN8rp/jMIPi8P4qNfpYEVwyZN+ALKKuP0Vp97w8eDrqoIpfrXX6t4CgF15Fv
PAoRP17bZAqJ35hc1CihYBmf7Blc7vuE+qBIBnt/2Jy+QW+RnNYvO54D48t4cfUGSsdKeR3M7Z89
A9lnlRsotHfF0n1hu1pKjB4VzhRdW7H1qHgcJWLoGCskp0JRrLPc6YRY8LY/JnhxTQj40EO9Q8C4
wiwjLBYyUGj81+9VB5eo/xI3gVwJo96ZFhdb/BybnZFM7BWuowoEro7Qd/WPhlConL3y353lnJQ2
xZTtFVuq9mgDZVjF8dfJgQyjg8ftlWxjATTLwtXSm9Fb9yKPelGjZXLNmuSbEYacUz/RedRx2vue
jYTbL670no3Hc77pMB7wcdJbndFzSynXIWnxy+Rwn/u22O/LDVezowIl+qNBUvZB2JhsJchjmhzs
yA6zuUiW2eSGkf0u3ywA080oCXMuDNXxet1yakrSwwkQx/8xz+BCIMvSsXpKVETQowxi778AYGk9
3UzzTnvKLuW5bZe+qK793bYND+WOWt3Uw0oBeo1d+f54P2EwgbZp1eAzLszG/d2EZczjTfxd6Pec
nNHLXL/kWuEDAZyDFIMT3IbkNH5L2dyxsT5oI42y1AhRsWAzyZ0E62tfCj8hBA/LSiyLZ0UK8eZZ
3IFKdULnZaRys046nLDnR3h89cfawPJUqbou7oB8UOo92U9Bj+1vEhhwBYNKQMPqn6Z2ET0LFw2r
tgiPrfCAJl8vMu3bUaUoUrnnodK0wBAvY5FiBLs26Onb3G5gVCzvGELVBr/kNzDhbl5FwBEfpMnI
mpNBZUEIBAOqA5ooyy7PdZPQmCE9pkIqj03IE+wC+aVf6948uFXaUBZY0FM0TsL3QlNpzDTu2Poc
sZgf/KkJrpyBb3p8kYmoo+FjIM6aEvwaqqAse4CMXMgndP4x0IGdOFkJ6eiv8DtarXOyUZWeIyus
w7BvL5sKa4BUyqbn/rLgCAyzHZSXtJoSBSgpmvvQOmjYryOYMMYiyOdwWkioqHy3NWXsMbX51R+W
lGRESUjksQ6R+WQ1qEtPbyf6FiHKY6P9wEwOSDVlK9/gireK44SNUXYxgWhlQODk7QkjIsuZM72O
kuG9rfLeijum8CHE2JvE0y5RUj/PO16QSxdIEaLBpq5cV8BMeSlt+m0rNoPVdeE4FJdqL1rPk2Os
HlQS9GDVJb4QRF3frXC9ISjmTRZhrWidiQkrG6CQA5NsBkXkHS/WYlhaOzM0ul1xpURsApzqB8nc
Peh4gtbDPIawRe1pn65cTnesyKmGODvTfnFLnMQHLThF63DygxgdaukaItO6xMAa+txhoZ9UiL86
ChI/vVDv6elbL0p0uLsQhwtzzOkrJrceifnvuzfHLZ80IwNXylAMzd8WPRwBIBC2bLeQpX/kdC98
BfIRmoWxh6EaH2OsdrtF3QMHbIMtu9xuUktQhUI7iCmjRaJvg28RCtYBHqaOR0x5PNcbKDMyvl0O
UMyZzvJJCP1FltQrm+RhsDuW2QRelBX90B7UDmF/uFbD3A+YAcyKU8yHtQEvEtO1x92G40rt4unI
mUSHV8kqd72GDBWU5WGFaZIde1S1PUnAwFWJIPUgttdaAeI3HzSNpiFgAs3i88KjQ3oIgyYefHq4
RxnW3ERcvXfIP2G8rnoE27Ym6CAfdG+hwML5gd2+Mgu4bQDWYzgY6ow31f/GwB5FYYdBKwR1T7Q2
/VK4PzvoLZ2tCRyYBzUbW0Lv3AOoLlX/Fes0BmQxMcg07Pm4E9UACxtluWJVs3pDr8Zm1ouVV0bu
iyKeWsNH17+EkKSE0JrkQkNcGZTdUZseKqOGIEDBsvBTE4gqhz1v0F/cG/gFBuJG+97buKZnBaDv
ScXEtF27DmCm81CgneJhblHMKee/XpugvkeMJooKuMUuw51srD65bshEbNfm/dbiw76fttYhoSWX
lO0dSaxLZTJZUgorWr3pyLoHnofcQ1D+JLVOAbVo7ckDSIAXu9nl0tz7rcht/RYAripVOCoKQuj3
4GoC0P4eGEmbiDh/s/K7/nz6hntMDnTwtWMPhfvNRUziPD+vTRV1DZrswjkZQjxflibmq0QPgxnt
XNmudOX5imvyx19YzAF22JzoUu3RDespzWOHHzI9AYacHQ9hXYgkqp3UVZzxAKWcxs/ao9toXIkK
wz/vY0o1gOBnL+ds5FGpxvRvfECI0zyzkEesvCV3JJx1ZXWzxK9BSVPZjQrZjrt7ofXFsyO3+fIu
iO0RgOHgT6HBRO7MqeHLAXqaZW1fINxQ2kuuzt5Gs0PXOJrflnXeBsD1fFwaMhL5dQmfkATqg+sc
D8TJ3uNPIFiY0XHWwTT1PcRNclbqNnrNdoNL2QukaXRPyhzhOAGb9fJD58HJVphstHfEC18ot10n
JEen+yIxyA4u+3xI0rJaZQwKYlyN6oRhiPsXX8HTWJByi5MWEPJqp42xTv2zJ4UzQe12Vmql90lU
Ghw11BShJ98+dr1CvTtX4Erbkd7hmNCB07PpN8D0oesnTyZGtkRIdrfa/F89qhXcv4p4EW8/w66S
0LBX0mDyKuv9mtWTiTxN302URtYMGA5TMXftRBdoSaRac6nZQUY1IH49TnBa9/taEmJz1TQf56xJ
5K94VWAhU3V1Hy7ALPkqeDMNIKK9xgvDSQMLsxSaf+Gs5sSJfUHGV3wh4dIJKxXh9qMTE5zN4pRS
ApLm9XkjBjhkqBI8lgMHnEvAAK0fFU3ZRi5URf3jL9n+/NoYCv56yxp2fdzPIWzIlniokD6+HpEU
OQBb0cTmisPdCLVE2MRqpPx9+w1g031bEwGsYdVlnDqMN9ZNML3EBlpf4JARY0pQQIQxCs0/BqED
v0JnhPKRm9Rr42a/BqNK+R026z/j2oqyzxlS+a2KNpb098zKT9C9GFA0jxStCltuU9suQz7bMQlL
uUQE0lAwkABFW4yQePBr9jd9JiY0P43gLddHXJkaVxZYf96fww82HwnAWS0TfzR1SU8gpxKff3x7
U4pW4hZ8rAtrR9K+TqO8vI7Fz3Fhj2UHA3fBYXd0chFo+DOp2KxB/rSeQV/7EAQ0fWeeDj65fMiB
0BvFnz7JwjrBB6sMWeiEeVW0R6ph8NEghCvDCkfqVYXR6VNszB9KraNj6hTLMWT9S2lQY6PcifoA
J8UzVnkdkFG/qjMe9qXFKjc6d0wPCSMMB8GtM0AOe7JGed2z6/+r0VuNSNYJnXDTkc6MfUyC8+NZ
SQuOW3fYov5EaSC+vaBYxLfWCrDpZvouae20Up8mJdy57FDrOQKamUjaldf2FtR42MOUkNZ2Vnvr
JDPAly18a4CjTMME8cZNVlA8whDEBttJ5RMsgZ4Bv49YxeNU5i4VJJnOFFi2o6rIKWHKEbgFXAMP
n6LA3NHQER1HvxA6NRL0QblYqLf4EQNeDuKA/v4nnAMuAFWSNZhZLRe6obpGhCqJmoPCC9XTA6lo
Z8J1dCqex1w1nVYgeWWWmBpAuiqP3gwaB31cK/440m7QZqjMO5ykkWPsZDRRXafShwIPBOQ5rC8h
ByBHS85fo33QRQVhb95uYdzNwEyharaOkgjo0RzU+KKzZKBqT7wfj47lmDvLqeN5hSgOHlbiLkpp
bTBu1P/PcgB5WvtsBzg4IiKw/pY1b1szuyBQytlriG95fUa3auIOJp+6JRBwxOeA4yKMELoSx1HB
lL1PlhZnQWA35BCsUw9c26qQKtufwFRJdIUwpR4fbuTvoNTi+1lr9NUsyhNOz7PlRscHbrtopm7n
jyFT7hkWuiT3KPqvkkpxkXO/fa6rkXnJGbDoRlLz6LBg+vXC6Uzsv+OAZba6c2cm72IkrDHtm7PR
ZJ96Z+xZ0/hjsimTT4wzYPRmiXehiLfMerfYHdv7dLiBpymwRkDNq+qQfF7dlNjI7WHAFEwhHku8
yXqhbTkCHCfBmP1bkSaRNaL9Yh/pS4NbfD0Kq3Ae+G/6JTLkv38dnsmy9eKGx9KLmPFfYLX+GqG8
pFjHtO/9SXG6COFdP7x7F86sVQr5b6Pq4uy34xq7F/03j6isRd/XRhaaV26bFsNpNMNnMFsO07QS
xRTT+QDDSOEB64AfpWk/faJNt9RJKHrENvLciyGGYierO5ZF2gYDv1OEZOlTQ02XZAs73q/OJn89
lbGHCoZiqmPD0nE56UXD4b2bryU+wteFDDtvLA4Y5cakSO6o76bIiLNODU7deRcBynewjtYUHKvW
ep29L7/GTJV2TlFVdA56a1qygwjFnDZcvM532PBGgkv0xSLc1NIVo+2g/8KPyZ97G0f8UphI7ECK
6odN81kFdLMlWvpHQ8YTC5v2yplr6HB1YPiUK20U3XlVA1C+LCPh1A8WuXwrmnMTd5jc93B8ZQRo
eLeS9surMtzvLmnuMFu+mOl4VZuVyXLlXBjVYk9HRO7Uj5ExeRd1QxJH5mkPDR+1kxNeAuDCnQRQ
bTbD4ZNzaZhjJWPFGz0ytq8wzWMsKtJjR08XN5sAVzMrcmZ96ZnJRiJDNEmq1i+7z2bjamyTpx3h
X7vpiSRMrhUcdaIMvbF07oA8ZJhb1pMHmpU8XEVh0v3dqyeB2yw1GLgv2WAa8QuFTfLeKgP/3ON7
Led3GtgeHvlpXrL18lLynLjoBN0OqXY7YHvM+en6XtEYHkn529TCuJcUiDBLb323rwxQX0NSR1rg
bPm8oXnAewaIDpvDhZ7awHUqONBWnM+iSVPw0BdPIcfzgbNvnuMOqstjCCddw6F8RnOR1aCZZsa7
zbVJmx1B81wz5wPWTgeg8q8QodnQGted/SEHFUQmRDX4ZoPBke/816ZoVrS7a6EJQvSv1gCR6hy3
WeyVBIjziZxU02KskWFamXo8ChXqxLd41wOHrXHPP3GBGyzZ9WRWdeBWqrppD4L6n1nGf3sm6d+t
v2k6ON+uEzf/Z/eV+X0ti7iNqd+yoiklgdHbTcdm8B4+R1+UUNrN4yXKf3lKbJqwGsc8zXPz89HE
8dXiM66tJHzTkCYYVdNhzYGxctiyFp4THHh3wJ5CGtsxqvQIjGc9frh6jS25qSJpnLEdh99yPt62
H8cX84Kf7InGXETI6btv9ZASs5Umc3wcNctyKk1gaHT29m4Z/2Bd0M2caU35Lsn0xAaJ3GddjPJW
macYfckWf+qTJpCYxfMCM/FtKvfhGiT4Sln++YVU00BdHjdhCBfNSEbMcyAI+roRBwc+L1lBZlwO
EVUKD35ZjBveB8Ff3Q3e/veepjg21RaFPZUI0VDt4u3uNPLk2A8NGTSk8ZuXUGoWne10g+j4D+HN
djtpBdMUDgMwd606Wv99gSOHCTy/hxQxWKT/Qgx45VnjPHzngOqIvx8N7IMyV2PxjQ7kDsYyQw/u
/7asI8Iayx9KDnmx7U/+b3cfoIhNHAobBHM5KWZdfgHbdtnIPhKybXZrGOc5qcbfH3Ob3mpPsDE6
A0nA5BK7GZxWIOVkO7ED/yfjrAzUdE3pW8AZnFKTZTNnqNHJGClZBHODjY/617hEjs5RgSoRpqHl
jiAH6ZZqYHotxzFR5RbPdugHzYuvR5nvaJoxWVZKDo6TvEWQRHkxDJBMFkVsX7jtwe5GhoiykBCN
Ig5+UdVoO9bKULdYLK7Pf/Ltz+EWpYQ8Zgnh+nhVtRMnYthHzlF2P3IjR4Pl8cTkBZ/dO1IAdhI/
AVYPm4QwqHsnXwL30BdbZcTGU+sfPSEsPPZezpmpg9Uf/73TyAdvkNwrk4sQP0eP8VKbXjWn+Cjx
Bl6AQdtpVnPrnmi2zd1hBdsHrINGaaHJCbHwgNPqYwJJkkVeN4P1UXhOg8CC7bx7oSmeahHbZ1Is
bR+2zt/KkIfkjlD7CZBA/2lBRhByE4Bi1Usn/0NDvsvWN5+WoH/A9oBXoSL8ERrIemvACN7Lb4Cn
/iecAdQdKj5VYBFXhx1iJL5vaq5PjMEgUbHRvMh5N0egtc/drIucNOcZIh4/dT+06CC/+oMO60UY
swE9V20CCUZg4EBK7OntRyaXh8kEz+uqlowXKZK4NoLa9gQzolRSj0NiXll4mXeRqTNXGWCit45s
VA6c1Wf244wd0/P7cBJZLxi5u5OQaS/4lTDMcddkdm1gtDIIrvLpWMBl7w0UBNzqnXKP5Cnn77mr
Xlmb7BYSgN4DO3NLH9htxJT2/YgCSWiSyOb0U1Ea7bx3vd25Czg2z+CYLRDKBSny0xCHmtK4Q3VV
jyb4vg0Vd8CJqTWOVWSxFdxRSt/f/e7tbPQTJcZUxar5hWBajq9jBpcAl6/y+nSL2DVXVcbLzKhk
O752sCwYVh8p8Hn02D6Jyj2nBE9MbnLRUyKEBuifD5Ng6boa98dBQUueD4pCcyElKBqJ2v9owwhf
Pq7ozr0v/B8mgSs26ji/Jjf1GOF7BMZjOmErfYdP5XiwJ+AdJKK7E23ErYSbqCMrTrYQlrSq3+Ve
HXjwcXsM0fpEVeY5AFc8M3h0F1+SIcjLBZXyWKr+B492PVJETDX2prrMXao8gDPvd+SItT/nqGyJ
0iVVdIrr+Kx9S/LJKr0kiLy8JjEYjFtI36OdzNztJRIgp/lxMVXF6M4BBu0lopTKSfS7zFBH3JmO
/cIURl9UBDu/qZ6TmHcQxrSoGW3H2PyG9uLlbjwPj0NWp/3sM/P6jTiLcMKB7FnJaDKfmZ35xEzg
r59cNbMZf9qcCnLEnJ9OTa3ALuiu0vHiIHTzz2cvH7H0laWZAl8IDfRgf+L9QC3TxToQGyxZ1ck1
gshTlUvabaZgbQAkRFlLmzO3Ev8KWEf+U0r75XKFwyUt5mjy4wZ9FGfvngXkG4IWzQW76YhHx7gQ
OppFE+1XZGADbDcW0aIT2bBXm9IJRMsJkivP/y2LErd9fFO2jOI9+mwvdJMm7c+93KXs1bcKgdXU
53t8WJcdLqZ8XhUNQBPNUfv2pvRG/cnSOKgXI4B9bYgxuhDBEjo4RbQtQ+iSxrIMNDU3HiKu6NTt
XccXvTO7ZkDluQnrPRHHXythIbshkPC1Ho4p/9n0cDzlJ6M696WjS4DjkV4R/dVnE7ntu2G6/ONg
GhgQXC8wtIxhXw3q79ZIdYLBEMyZSKQ+XZcKAZiZ4BE+/ZDIueSPedV6heoIUrncMyk/e9skY0dP
Z1d/Cek95/OaEhfcMyhiDQcBXLpmGpqANnofB++7OwUJP2joIfirQGultO+/0WfcBfd7Aq8g6WyT
OnfMRCVLlEXcjdutNcUCTlGGfKUnnUaKUrZI4wgpLJpK2K40IvxiXXvftcakunl8t/xly2F5Kuxy
ZZcyD7PlkNBxeMdDp3/yqYYs4nRnXHXAvO85FFbc9T10AJ0x6uLI6snrLxutf7JiW5jAIOZ447Kn
NT6ZGbI1rBET7Fhq2WdRA+flpUMRLNyxMrDuacTrRTu9Hyk9W42GTAjIRSofEX0edcKYre0+VwDx
XGEc52mNHodFUXUtKF9OGtdTZtmXlbG8CtefoD+G+korrxNlt1gaN6dbWduweFDMvMrFWD4wxvMF
LKpwIL0p+NBp9tqj7xkpjNTniAL5L+F/+ADgbBRpu2oYAGayzi3L+kMP3nxiKvY5eyY8h4qWlLMf
kaVys525ZF/2He//0hAIi8fpV0Z2oMtxskrCRxVJ1IGp+DdV/WTojvWogjTYyQmqALJBIYJv1Nrl
EYA5UU4bcig7gRZi+Kxz+GBUcY+c1SUgvyuxHF9/ZRWTkS37+4/3RQSiH6MdJJIIG5kJ16WC5wGA
mGfWFbxwzHlSjwIqsxtn/MIMXksW7coutpQJ6OxGlHfUDbDdfz/RTVKmBhqP53wxwOzAzHwQ2vbH
VTVf1ZzUyMqquOgJDXThyxEFKS9x7CARNTRf5XtnFv/thBDHzNfmSstZL3d/SmUhSCOzvnMCEQhI
CDR/WdRd0fRiigp4sTnb7blKZQZD+UNrmZ0xW+wGbtByTn3uvTJk8XyfOk8r3VHRZwyhAbpsSls5
vI/pm1Qr7LuVapX8EkRlh0dwdnBDMAjSb3c9aPBRLFWB2OMHH2/RNAwTulwfwZBA5fEaBfXp95uU
2u6LjvT817PmAmZt4xdzFzBVvuHYQcUKXyMVhCy+XdInnBYn3RP5I72t+pyFDawOa2sCA57UOxOP
XppXIJv1N2T72gUHY/QE4JuaYJsHV2MC5um91vjiof3jKraLa6Q5FfTk/daq3YjMI1oEJdJNMNFG
4jMaCkUpFD20/JhYWoibrSE6NHzY7Eo3fBWNfivUxVGdaYNZKOi6lfSReLqixQMjxN9oMaAAJX4z
Anm0/KTwRXA8udNL3j6+fhuTJrTvnXcNYb/pKMqLXurq6HVYueZEgYWA/lTJFdNJOnoHrsYqnZqN
EgnMQeg6yFNVGdz6tXqiskma2KQASr3iX9KoFQprzIqeir84Mn3aIS5lEYK+mg0OCrgqd0MUSijH
1OOXgBo+Gja62GGCKPwlYz8nnupvc9uO1iohc3BagL8iwbrOudOEcTsVw2rjk4591yoyFarJcyRx
V62bLj3kmbDEcGXxUGg/VWM4LUzmvUjXS20mu0wBncJGGFjn3R1KkVQaFKRuoRDbJcFhDiDz7HOw
V55I0V0+bbc8Jvknw0+O4nUT4kFIy1fO7dKYGYuaVf+q7zGPUVnf4ngJK5HjA6Mr//IMl/1Wi1aK
83jTeQjMhoIiKJK1fRXJ9Su+O6lX23QJCeMpwwqbyko0Zr+CUKU4wcWCFuoq8JcPyFes7Lx5Q3ca
trhN0q1Q0mhE2J3GmH/hcqabb+QAfxcjI0ei3PHSxWXtnJCwdOYuRjl7VegG/XKWHwXDAc2oW2UO
K81MCOTnAxTnSYj8MvjR//VFcJ4UmFla6z2plBM0vc8vJ8KEcVSx1nzPgOx1V8kdeqh3OUqhet5e
iPLtbWXcickOZ+mxm7Eujq25WZgAKAl23e/do96ErlOf7hiH5Frm9C/IWz5Fo2wj4vWEoqVd3MZN
vBrrm6IS7v7AX68iY5hht7uut8fl49L04G2FW1mf2SulT99FGgDvEt90UG9vYx3OdOZWiNvaXC1/
HQNK6oTd00lBTxkzeyiIVxsA2/fuqADeYuKwSXPLdorNpuSPtNm8qTLqGhY3e+E+20F4ccvSx+IU
UKBp4nmaFR12jtn6ziHoX9ujcxl0l3kCjJjnw+7dLuPZPd15aKCzTWpzqAODiXyF1Ku5l7G2f062
U7yhnF8v8WtJaB3TNqstB5cmE+Wh3FnQSCUERDSqJjulTFRtdJ+DjUE5wOhTJZzfZg44xjC4ODYK
UDHcbqsIWWQ4QZ+0p4AxK9PC8PXGG4pEPvx3niPpNe4e2WUPcTUoR7BapgjFSY25KWAfANvZUG4/
V5/2o7vIBXMyw0Ijb+v8c8vZWen/0SLIUw6N1oKR23j2ICzU7RwAdFh5ZIVxKadz8Oqv3X9FhgIx
aVBo4h2q4b6VaQgYTepHY2H2j49ueId6jOa7nqD903XX6+UbV6AZ0rCesAmWfAZWYLO7Mn5Fb2tw
lkoVnBLWtY7Hy0zXPphNO/PXFemlZTrTvAeXxNMvXj9rl4oTpzoCgyepjZQeeVZDGYr5f4I753Hp
snAZUdL1pzdjpmfHSA0MbpgrU01nQIjvY3jW5X8dfrGykdpNQSxFD18JRp6amIQLayz/PIT2wZco
W8lY1RiwY/eDswx78zZ5j6bfUbr80yHEsDjd/bYkRTioS1Vbgzi/Bz+wVPDxWbrBChSDcSf/q4K/
KLYA3yn58Z4ZIvqiBMRxGKCTfheZ+GXEf2cP/iadJWh30ttecxL5UNp+Pklld43j10HJJRr1OBK4
IEvs6Qjvw6BpPutxlr085UdiWzalDrypxgnSVdE7gkueStpDRxaXjTWgicv0o+d/j+/b9gDMo7is
rttB2ohGj4OBuQw3IMU0+6zN/hwyBFAxLsGkehRd150l9n9x+wOGaOVcrVn7cFOm0cdd8Z574Jvr
U3Swc4l9QHLkB3tsVtVu/5LXBWrk2vrhqxiXrIZo4E3r+CO0EZDeYrWypDw4d1kHKA+Khakmebmg
W6kq+KP0oReOmcXiBJ0XE7SBjgEmJC4vBM1wF96jBSo8XSAsyAY29/qK2mfzmpMXUfs9/DfcIiq8
6V56OOuL40bjarzmRxrm643X3xquag9CQJ3y1bYJK1/R7r/eCPrtrGJZqxNBf+XjTPtAPcfhOb7R
w9dMr8xOxQUVweBcChtp3myvPcjZUSiiP8VFkFlMLptfyMSn0SYgqpRJVkhP++m3sVFxwiHQAwDe
bRmBLz1EjMm8mEaYsLJovI3tewa/XM5MpEkRB43VhWxgxwLmHMcs5rogl5BY2QUIeTqloNZSndau
moHk165OOPCpRHd8b8LmH1SAy8dRJ9x2rEVpzKy6l72FR84UIGWEwwgm01h+WQ0Hc67+lRpbx+us
PTLdm/ChKcAY38rK0CnMlsc/WT1q7PW0MQB8XLS1KQr3y85RhaVrhJntAsEcvgw08cRUPxA/NKBe
IOI2UAXBtwZbtxBZ5ABmEwb7UsBQSUFjNloEc4uqX6o/ipm2IZ2ns/bwqarvMkw4IXbPIDQgwbGb
U1LVQdC252HfezIaiGXp2EJTlRGRAqkKoRD04HGDC+uhDs8A1Ezbt7BLXciBYx0T6AUahXon+x1F
SPxCFrkqJ7iKgNvILqRH6toWBj6G5Sy/LBzR6wP69UuXHr9oNlQFqao5aQ1nUS8UPU7XlrdtTBPf
ZGVpdZI9iEgXQlzb5W5Kmfj6SyRCkrADmD2KUUuqwho4bqFlkyh2EtY3fo6PQoMa1MgyhZk4+hsW
51tOSsJIkBxEsBYtKCUOgWc1GLbGAJkXX7lNxR6/nXOQ23ZHDaj/mz8RaaFe6DrBPLjHXGJP/xNS
uze1jZIdAq+ZRekE+GyF+ut4zmgVTTHAuDIdKOSlPs2zPti91xnThMlPREA/kUbM6mPISvT6FSKi
638VXjsxjQp6t/ZDCWXnEO2w3+d1fAu3ZauAQYMquCj2HqGbrnGZZT6QtEH2oNV7fduYUcWkATlm
ioG+N6Ik9pyuEEkVkVRoRbLvYWG+faMXkTH5QGuDcUSaiKY6B3Y+Z03s5DgVT9jUlHgQo0wCCJEl
7ubnp89HuGNfM0+Lqg9OJsWuIsrLNf0thF3IEuLdqz3qcff6DGe87xGCmwDlmCep2QzSJcuu32LT
tpFAiNi7zLwHpMpt7hvWhy44YH5nj9IaMbJGONo0LlKj1TCP2OXjxuHiVra97rGqXJQhrNgdQE5Q
ty9EnmX89f4ytC2CoB20imC1dUdFLnpPXIg0YU5DNkLtuo8kSEdQqRuKpWeDHEmtI84D967crDG5
asbKwQxVmhEW/LBLFoY1tyHxu4+Yba0Q3JaKW+ma+CBXp7oPGaLx3sBj8IkV/Wsjme4WG1gEsZP5
CrMUnRK0A1WInSBFxF6zgjvVnBiRoLj+25JkRgYmmNOjx+ImdWaVMeBdBSExIC2D6E/V6O5quPJZ
uSOuUo5jtXfhDN3n03+tnGNm8Qquhqh6hXlG+Eoys+A3Iwv4aXTJ4SWsx8UTbX9MbErJFtjGqsoW
Rj36lc4fxXGlMN+uSA/aR1uBCsjPe+uqxug8hdiWgaxAhwwJndY6Qsd/ovFaF+N8WzB8UM+c+JEF
PddRvK4pFzyq0q+gLNe3R4gx4bJuF3DKUYL8JHIuqm+r6syxQPI+D/HS5TzCCOqWsmyQ1HcZlEek
OP7xcHg9B2Ayg1quYVdw3Ozt1VVWPNZhI4Ez6W2Fkzinvzfuv/pLiQg/IQFETqyB1bnd/0Kc22Sa
dxDpVeKnrltAugR8DDzfnVSF66CiqUfTlFQOs9cK1dQhVdub3ZLSLuStc3rcpqCsnqDHRhqS/Qoi
Gl8Wa80nPj/vunWjRXGZLoPfI9mpCF/zut4d6bMhJQW5uxf0uSpGgOyKkeSNzIDmYfnvC7ZiVR0v
373r3ja9tdqGb5ve6HqpySJwMmgauqZzudfFxUydoHYfVL2Qjlv26O1HKR6UCizsAfUe8wt2jSe5
C/nyZvsjmtuk5GmjhrgjJExz9h3VjaFcqWBkZMvFhDClLZwxzSEwXyFf7lA2TfDYrP9f1TYqtJCg
DPLFj536mes86CCsbocQTV6u/ab5zEz18HYvfeCoDF/Y3xPfeOJcVzTrtDdkZ/2y1uyCU6QuasGq
gpvKsTRDdmHgYKBR1zRZNR0vBSlGP1y7T9QoJqO65jQNcGwyZvv5aG6ee4TvOQwFE8n2QDTruFfe
G2uG/CyilFJVk4xhKG+8m0JoHU/6Tbl7ja4O14Fvk7jC7enx9jIa8d24Hub6h+RHcF0iCxUIYQW2
tm+1DkEZVnJQSSazJGPtL0n4ix70LPeunT5iYvN0fpiRhRMwmnBc3Oyxu9xdsIFRo2RsV46AC669
uL5OdoTXuJDNPgh36wV/Gfshx8OBdAPD9djrfNQGkVhXBi3gbbgnI6NHin1cYB+io9EuK6nOWzti
8d1cKartDoc99QKh70Bt8c1/zjZ6F+nhC3EqcObXCHbffDhyCQaf+33ga/i7vp3DAAI7URQKEZY8
e9NnyRJA1mzoJDla8EC0Fmo34G0ER+LcS1IFI2koQ7RF/GUMcQoPgHzCEWATh6f2qlgo/zqkh89m
tibs/loM8lGG/AUrEEODDcZzPKkMUVicflFBjGZp45QNHN8u4ZOZ3BxF9T3jWOww5ZKv3KQ5sGty
VCF/ZfjTGKH6wUoV+3hcP3wlWrh+TAadOTmYzK9K5WpFER6zVOxyPvS9rlV+qf4sBeGfkpfNIPTH
Iu67vEpiJcexSap3HEq0LiiZrKIJi+v6e2wl5iMXzGZX4yk8PuoK/b5mC2zpyVWQDHnWxNDHUUoR
Y7hgEF9NzVbG9YKqrPDqpAx/Kos+Z5DWj3d5Nh5BRoERaKufykLalTRn7tRudaD4x7+cfai1Cmi0
qTr5ULOQzZhfIBF9FtB2Qnb97EtlY/xjgS1+IDZggcw0+VH9ucyoJ3wr2qxvukKlJTwFVRCRI18s
ig8k4WVM610nsI6DZzwcH8ALMJ1dYkdvZjhrMW2CWoMyD2LFBwvA4H9OT9mZgRIuh10bOO1rrZad
oAvPaNwvdm/z2sFKbW4IBrEmeRq3zAwF3XVtfxlCvC2Egfr65tQRsjDLzjpBLNGNucQezFspenHV
cyHEGPIVahXv0o/L7RLlvjmCPiCADSWaVyIPYvDKcOG0mz5nsplRfC1emmaa+iiqKxtELx25miSn
HcL/YjEoRtNq9MXsoweUCKADK8AvNEvj+fTb5+UO0f+4+S8l4YtBTN40ThlmxMksjOv2CUWqKUZI
Ecbrbl09hpiajEv4IEfhYcvaNn/eek5H6Honw1hXBrBU3ouja+ISHhXcpxXHtu5wtD185fbQGsXj
DnlejbQzco6WVTjBlNmI0UD4HUE+2HnWq6NtCHl8KCGnHCfNB9McnzUjtPACg6deWN7yCxQnkADT
kSoM2GhB7EV6fm28/BBAplOmXm7qpzsBm0b+Wmh+kVXN4j4tp09CjQw1EYRpxdob2DfxHSBGph9Z
tk4QYGKKUXa1R/bYXLlk6sP61AiLYQPXz5ifR73suFsa1o3iS8EA4miWnMlK7e6f7l1wj6GkNkuc
g74IY/EPFcl2DL8mt7whuIA4mHixE+xQe9gYlcj/iLz0kJNCdfDOXZcDepZSY8PeUAQTPOMh7ADg
TEi39feUf4lb4fREJtvJMcAw6KSlVgMm6KZBSky8fUlkFoZRm9Svp8cavZ5WPEDcdRrSk+UxPtCb
HxY1tg5OkMt6owfdMusfHrk5rLQ+lan+yi25+ckagDR3rlMdAGyPpjNxZ58X4vBDm71J1mKk2iXt
VM+pAsMxtOXebA+fTSXfnU3AyXgSOkjJgIKmBk+TBd3U631XRi9Wm4pvifmeqA/IoYjss1MYCwgt
9R8jEGyrEoHW9bppORouJub7WPfYlSIhBrlUp5g6zYhkQTCWNqO5NBZLtUqQMZeXExMLxHundSNy
bg0AiCV612xCbVOUoqO0eZ+ZU/ns4570OD2PFH23/fVUGg6NZxmHk0FLU7RgUoPMvfYcrs1GTIsZ
oek3ly11ZVxmGd5pMLA3MXXECg80LiFU5O9uyZGDlWv0R5OWGWHQijjt4geQMW6yqiaVDglzOfGl
uWHJKWnpeD7L8YItELbIuhIseqvorPpJf/Hcu0O4YaAO1dxJnEEEHAm5OQSw7KfSE0dt8u19T2LJ
9Bc7ubgB+I/fg4VoaXHVaV3vyC6gAFd5D3sCatHJycAQX4lKoB5VNc9u6smAKzDDzpQI7xR3dwss
MrwdJhj6KgeBHywY95IvepGze+DK7yc+Jum2Qt0YmhFPGk2jNC0DHOyO+69b96/cPuL/MPZWFV8c
nZt2FK1uN/mlWYjNC7ygeCW0QD9yj/fTQ+StePt0b+gdASZq6MqzoBJ0S6fnvajCC1wKbAvs2P8b
ZDzTI+3WLEF95w4sOLkuFCaRLfoyxHQzc70Y9UxU2eDAUYu9MLVv+h79pENeQv2U7wbNz3rGhcH7
GtDSDjTmUlmGa49ccaoY53Ss5x1GITtqVFVwa/nvkCiDgt901MKIoSj7VW8EsY8cO09SiNAPhfhP
37ckNICvlM6lJm8JgnOa6U+1YdCdYS7DJOCLqBoiOIInn3HiyIIVOocTGSDY2TvyRIRHK2g/D4ED
iIy0pieFBqRBpyFU8Z8Q9SZRdocTLH+aCaar19Eacu3sqN37/aCJHn2awkCVBfc/6mIAiuw9twvS
7jtqsPs21fV53VI4yyhaXb33BPRcni28eyRyli5mJe1f352+KKhdBn4mom8FiRnRBZBjltDTfwyE
Gvf18fCd3HkHbw14ewGw/lzu5ipNhzGeHSxRld88Nb52FQzOJRrSGxh8zCzuUM0tUl/Sbcyd2tox
+efquBvEBE1AzifOWjkRb6wr1dXGKWRUhC3ovdb1Leb2FswB5idABeA6DlyEVrpj+0OFP1zM0v7D
K+Jdndu5QC8FbnSf+++cXgDl26Ji7mWwEJ5nLlEUAWe28So9Dw2BU6/iAguOxVEiVGvvwncIIiGj
MO8T3GFGPjxq7p/P6NurOlYy4ndETb7NwrWOFiVel7Dgb0yQa8hD1sA+uivPqvdoc0jVqBf+Bw9n
ZPGaJCjXdQAIT6FkRQzkumIVn7gZEtdRdm0+XWIy7RoSNKjepEsllyMng7BPzYEEkDgezPXrPE94
66MvwqIO/15rhcmAxPkIrihw3DvDit1FedaCD14uMEIdEQ/GBJVJqdQoNhNYwpglBWJD4T6aI99M
ieUzyDNGIwXK7Sx6u7DDOmUurJHLPDzSZLfMJRRDI5HZNrPyV9OUZmgyY0tdopWyg8nmYHTTGvzT
jZbZgY7HqmoKjxtKORKcPQpPZmLMoHP8+YUkuPonURSIU692qmrNMmNT5Clc1PzMPua0ZeuM/HGn
Xvg3Zhl3YtgM9Y/KHYC8+O5/aYLDf+u7sGKzYExHbyHoDs8KDRLgEfyayDu2Y4GMLBd31G9KFPkn
hi7cLBrJ/YOuqRyLW7xevmH3JhWISVY0TbDG1VKpm+E+8HAsC5ZZMe0uqmq5O2t+7er10M+WYJxJ
A9LYWXpxTKU6YOrLA7oQyTmSHGox9zvPhaV+V9+zEbkzcST+w/vkdm0JVOUNl4lXzsfJQdqx/uzl
1IxSk1KA4x3QzSvzaw0Hj/49ujSAcmf8XgxLl/TuO4aH9gwwaFpRQMXVj9sq+WUHcRFvrnThX5q+
ZhvX4CoyL0l8F/tq+yOfZmHRD0NwKgDqxUnAEVE2urSuLPBo2AcYWSF3Uw95jl/7xjisYHPLPukR
cb58Bq2diiYbh5rvAPFWyIub2TPp1W/g7fvcRc7/FOOUKgAXAGAhHI5eexrkhEOlRQy1efV/2Pcy
hH1ZH1++mYqWf0kzvV+3/TuIsG7jPpqU9sToM/CG4oSVbicpplJWEU9GxhnXPqJiwccdkvJpBiK8
bHRbBPlXau/JSH5InS7gcTXNOPhtrQv1Iro9jXnB71J1KUBYbVD8iLU0FTRgZOpX1bLq+/mo+N8P
2jdlt067c0ZQnvGTySXx8GxZDTj0mHie4E38pq3su6Lf0tD0dUSo2LOPL+VZvgKxNscCvUCB6Gmq
OpJyRSZJ83eY0TdWXGIKkGfQFNFcEyLYBsJef0UtULuLu4gqjwKhVc9hFJQ2qow2woxJ8OJylPNL
8GV2STWIodRI7NSgBkPbRtSUnsGbpKe9Xi3oYZIUW76fhiSng+DFhQyXpqfNmcrMOw6DfevYnHHE
lu+Bk/DyX7ihpWtXrjs993uUSTFoWsk1SwydisMPsSTr0TU1Jp3WE717tiEfyifcOGgew+QzCwOq
jwtVb3apHrokNThqw/x6MSgIp42gGR/xnGsAOEsO7m804YaFZZv4UDbcdJ9kxsHP0k/ArwRgSGFo
kt7ZyuPClkJcxNlxHOg8VskLkblPC4sGZ77oOREoLu1d6OdQ2ItZhDoKkzh/MyM2QnTZxPCSB8CC
Ey2SRsFboCC6bY8yU/mwgB2KFf0agKdrbSCAkAeT+en5YCl3/RaBkaRIkoP2VHLodgl6YlQ7OcQE
jPZoTwq1+b2MrBwjaL+h/L0XgHnXvFG76Jsd7LOZC73uWDWQreX/f7sgleJS2VvfHLy9Zod3t+xd
/QrpMMNyyUeN1CAhpCqI8ewEZrC+1+diR3ouHa2MkxNT3cX22QXC8njtuPfbj9Xh3EFUgXUN/sTU
Mml9k/c9DN4LOVwV4SgdCKnJBOBZ4S0tWGbi83IFmxqLN9YzYr3kdIspwpo62UgmRO5TpEEzSYgR
+ZjflPFxqOHeH44sn05ncpf3X0LsblWUowbGwkjwC/PSUSoLzsV7uPznhFHSeMZsFl88uqH19EaR
ztpwpKS5FnT4qz3ou6ifXU26AnqnQEBZfGkAGbUVuiDY6MIbyZivvKrZ0juHrAyU5EREP7iAksfZ
VomViZbzCfRyyNmLatlgeSks3l5Vf6MSaID1g18cGTfZNUIqUrMCbSEk/n3pThV616K6vB1raskc
tS93jlI9G35qqZqKkweVR1Xs3h7jMK9aHj0ZT6701kAJP3Nbv2+Kp7xhtXBseS3smJpt4HyEbT2y
UcyOBIX6RrdpsOzBcchhW/RTw8Ny1o1XOuBzX1RAoNFlwBt/HAEyXheWIEXtQkT8S8Q64561zAA7
MsCU6CCzA28Qo08b9EzQxu1tXh24hRjDwruuc0hNPuuv6CdgdUblZjJEzaxwxtC513XPvhKCsr5q
cYPqHZtkOt8+j6iFzUcX30Y1jO2BDs2hmr//mfWs/V5gkNXCKCv06y23ejoa3UMT/ggmbXY/2UCv
2YBQlksOsMgwCV+Hg9RXz+7ED6EsA8glKEJZzUYIuaQDutg2yxuqoJQp0vIinQx6Rvnz3tqhSw/g
lLblvIJDVbj+6jn1HFlGI6M5CymLkxKXRgnCYrJxXv1b20UMLlrYNeTLeyT1nQzvYmfvMzarwKfl
n4KWEC6hKNnr4MzGrScQkVW0zLArPbRq7Z7VHbcnpKEItudKyZpI/W0rrmQEUV8cLtlbjcYNwbVh
OF/ue7TiGVmQDpc75ILhWRZ1w1nnw1cZYnE75ccFZlVjPL9gsp2vvS/P61n4/HopwHOTs/hsaYWG
93CEFlIEFMU666VYP7RyEVPl82j4ru2ZiCFmUmpJQb+sLCqgFpNG0mrmOMgdGAU3URh5EY1hnPHs
jVFGZAQSe4NWhkG+ZH+QlZmtYI8dtE/Ec+Kg9v8J8jDBIveG7nxUyGSryd43itPlqv8LBD4MbQ5T
DIC6AEDTNLXKH/6h8MCQj+rKf00bcwmNvEeIUM6am5OkXKNOy/mplMWkg4hjfWCLuwX7dZ4+Nl4e
HmIeQTKShJxIoMR3PHHjNHrkhWyHqEO+64fUWc/tTY4GA0KecsRSMNgY/F2BB48tefvI0btfjyQM
jpwxgh0lZ5aNb0G/uwGiCyWRaeuNJznbdkCwc8qWHszYZv8Y3NwL8J9LnCpdBXEDQ0o80MU5APFZ
X3PkizC1s8ipKcQzL57Vbk46kEpy87Opr0+Oc/att3fw9aldMBr1IxehT7GJkgnj63G2xS0sIxv4
x5+5K8iWmuNgGj1TwM+xqubm6fMvR8iV56OJT1/tqhRWYJDIZZ6oCkUxK/rYSS4Vqo77cewqD2uL
TBaLrPTDvn1V7TERAif+WZ0d4VzqCjqf61whvLNAGvIr1HndMHPnSfkYjYMNx/63bVhTJUjkzQ6C
beCR5jxz1tyNiPBwSzW27MObVPADVfT2WUbVL/lyoc5X3OWcidrtOQrYNdvj5yu/xZ0Mjo9GLR7T
M7XHTC0yjVMtXxsZhFLwkeDfzLbsx+dgy3vRwBTMmkgQ1tRvNd+RWlB+5kSIuWE5ZCpGepApX7J1
juhXSN3Xbv8hE6TBumaqwxpd1j01DHfAJVhJj4JFHr6m8darhD8YvQo/Gxke/jfOTFXod5TMPhZ2
Fxb/76ZLl4z4SrWqXSaE5b1u3G5K8wNgHC4DVnBs2FbI5+3AGVJrF/aiN+f18YcyA/e6ulDx/1ur
C0wL/cahoqYucfX8qGBUVwAah4bprkuCjVXu1GhK4P7tx6vX1jUcp7sEn68rdoghfl3T2wW6aB52
tQ5udPiAa2sVzFM8S+4Jsgo2B8BA8kHnGJwSYe1gQroOIhKe71ymolLed147LI4T1H8VwLPfyRCP
NbLtxJmKTZxKouYl29a2CDagg4NQpH/42WZuwkuid4NsbWUJbwzd84ruhH1a8TPqCO/6Sf/4Im2j
57CIIhq5PpI7xhbX1n29C3aaqkvvnWZGnx73tUPY6dpoeuVHpbhM9tTT919hFm1vWeey4xw+vyQ4
XivUmVhCwsNw3PPe7LU+jKyP7bA1aOUaUG3R7pxQU6IBJc4nQa9a+1SeKhef7BfBq5jGZbcfSgEH
kHtjvuxOyE1vssTWicLMeHaQe8g464zmUHX4RFip89pzqld3tX84Is+tLY2h8QukP5c1cei4o9ba
xHTojBtM/ozKEcGVt7UnUZUHxFV9XmSFayalWCSU3lEsgH2wcrAe5XQ2aLglLxJmHpZsfUvKA6/O
7U5XCtnW9P45cYrcfqrSm8mH6CNV65hzcsDBG62tmVootfwZ4VjxIlyfFZ4r088t1mOTUcmCPV22
oWwT+i72O8TOqqg3fvP6yrYWYDFkHLeXwNs7uOLHRyuyyOEXCIUAi77YlQIkGDT4iRrI7/m40eAb
93iJ7vVHV8dbvjbcq9ngKocerl1GcaKHaxy0UiBbghrHTJGrSPpbNXQ7Pworxky6M8rWOFpdjtrS
KmW/YH94IvRLDXvyWWosIpcuL49BDAUcKvjgP+RDsVxOwGZTlJgSPlJ15XpmA9Js82PNGyOL7QYp
7ckoWJQyS5sM6075RlGPZyeJsSh3RwFRRYh59ElDyqhNx7uqTMHRX9CUJkZU3aeockwRpblhw+zZ
3z+eqW6g9YCnCKA+a1tFpM4hPDJmKgpXA10V/GCNTMIfgOSpJLqUwz95B327DpmbYTnCabELmq7q
kxNa3uPpTWkCblOvwEudM6q/1TYzGxhJtFrTSc+FPM6Pbka5OXSTZrMsFXLh/E3WVt6I+Js/JLqd
j2c7dBrISUUg68XVOk/OFjhEa6kCZ3USZrpHQ2ZsCr8HmGtuLcIIbZ3YHX4Pe53LRDsoWDwp09bm
uBN1StXD+hPHLNyM6kv5Wb666XXvaIAvB+wEPV+/H6PQlPhBCAPxpuCNqFHKoRzxVMKjNdkF7ocA
OtY/Bb/jIOK3H+fHK64tGMCUh9nWMQsmrPQ3WqTqrxfMoSwEdDUbXfU7nLsNOGXXYRzNq5Oi21C7
MiNl9orsz8sHytlSyFavWsJhV3NKD2zPjfkpLY3Wa4arud0hj5zP9wXUjG2+0WXVfSeKB162HyYp
1twphmrGlulSygUYJBlsiAyuMl1n4xNB+9OKYbrFkikO1BicweK7z3NazAEn4qKtgH6Jhvwvqmx6
1En17g+K88dO0h6fzWAMLBmwpwRhfm1zsbtlVAxlFdq5ilJ7ZUjzZ4Zw6shv/KN5SqomWVEhIuXs
Iwy68gPLs5VJJnsm8bc1qRwXoD6xA2Fsi09GztDlQmgUxW2koBz4HmKE0yi1wDZ4zVNo0M8rzuYR
wIyAr3SUx8CSgSulIbwDYJQ/BxxYQ7aWDNZ7DyHxWiQn7sMP5Sx/r5Zh4SZd22v4ZnMNQmnB+uSW
7/O58Kg5g0nseIjN4OxxERxp8VbXFhBbF6NNF2Ds7aK1GWrrevUXxP3hvw0JyPZWg+90HS5sbfVf
3oBa0Ehmww1m7iO17akDWn0iq3TzNeX0pjW73qW0k7h5PBPKH8VhMCZDyMchJE3rsrvJDIxfc2+R
VfbjNwByjEuxqO/Ld4GgMTorGJew05hqRWPNa4by6nRqSUSRVAAOKR+g9KxinX64WcxwlXH8t2NS
xLmO5AUWwqF0AJsbbXxisIF8ptG7CoXibaw8apoBbP6jP/wVhDtybeEsMlu4U+Rk8Ph7e41/KTas
fZOCU5PENDnSnNo8zugHhOyhq44FSUCIWB7c0zHpRsDau3jWXPALNP7H81y+hvAuHza/raDoHpuI
wxON0gPHc3AN3COZXWKUoWyU1uThOmoJrIA5QOgp5aWFczD96H5vexAjhChngUz9Pjs5FYD1wJkI
7F6HjCSSlgi67y/kzDfciiWPMh21iV3Tu1jQRsQAU2vyeRwVj5PUEhroP36KhslSH3nKimUY6ROV
BBpq6zEitvosNFphQ/MDa6SOoKXoqnZ0K9JMLJllCB3Zgp7jdLkrb1sS+TRxmc6qaxaB1pK48OJF
9T4N4t0wSAE3A9ASOonu+eVdbwuLTatIUW66uej9t19jpdtX8QW2tcZ7SOX95wQJx0b2495H57rq
f+c1GeglecCDXEGnWMPjce3EDmCQ/OtLo8g4xXWiF/t8SoZi04a9zHPcE5MHNUyJYwxS+jDiNmJ6
morESAIS4sqyXRRGPj4nhejA/fbU4LVipX5XTfeqHI/5Wsq7RWIgjk6HWY9gMXwYMF+D3Pmd3o3W
ARc2UMkpjWdCboH0dawEbRyvoPw28twt2hhqwfQEc0gZWXVXFwZ1NV/QRwJS2H6PPCXCAtEBsEPo
Hy9fAu61rZGqXpsuqaj4kjQBmrMJkbxzGcBkWRVIlJX8HP5QE3GcJJL0Ac/iBkWGM6sdTMRFAIAx
XeGiLLroqW6H4pwu0DV0nXYYkGmiw+X1Czr5AoIQMLYTWNQlvYFteYjBmP/6FWkzvnuTW0pfmzgn
iuXlmkI0JGAM+2UdobOctP8t2yK4CPB7a4YdNPqEHuyFM1sU5p6n6YcP12afCSMfj9lhD+Ac6S3x
zijA2ZffRrER079/JZvfgCIYYnqW3neOpFBtEgaZxX/28VrCsFJEq4iJEV2HkjmNQUOLxHN95gZ+
6GZbIXVQNZApWX5Zh8/Q3Z8DGIoWwD75FitL4KqX5jC2Ekrh78VDMfVQ9ofaNNG31QIjkvdNQP5F
XCtBVKyRODw3oYU59Zmrr6eD7iWRpQK/gtnUY7Nkd/xUyXCyayM563BXK/UWj2V+EKeY8FWBFvXT
1vAD2cmuU/N07Xdt9cGBGTYS41fLYvhWI41lUeY0ClOB+5cHs6xKCnLn7rMO/L2iI5TmSHRKlumG
D8MnB05YPEpqSmEfq4/p68rZ0aEDvPfA81loRc5QkSEkwTuej/FyRC+63bE5m8azq0huR+rh49sE
KJJZYXNHWwsQjJscqa1V5ud2J2GQzoky4FFKiYbEBQW73RoEAE7fFJJed0PFopbsAkAOk6X/cBeW
rgwz+mOj88vkPKXk3Yk1e5mxIsELICR3Qiw3ZFloMDkxKMY1Z/cw6I05hWThaW7yn4nef5Q2Bny0
xd3nmJrLsQejmcG+Mf647y+iL/qA6NctGz584oWjQxM4njcUjoKOrhvd113gsc8g3FAnA9FLq4HD
Px9zHsnjPyFVEnyhUI3fD8DbJqXt9c1/rAPv42JFDTwJ7eJixlhy6TY0fECOw+kvSVC7ZYY8LMEL
TFVMbU7yK27ozHoKof3hgU7FirZb7jx/GiqoOIo6915wYzpI9D08pssMSLuZDXZkTOhxxotX9017
C4V+Q1OK24kp2GDUnmeJKX8Nmq8x8W3k2MNNyLUgxlxEvYDo5Cy5uYa+pb17da4qca/9brd85ekX
uBwpd0NULO9rACrkh4rlunS40fmxC2SVx4489Ps0od3wKhuftqaFRVhWgfTRZfROQEe/YC9ZdIiu
7Kd7y6IhtPqBbu8ol8uVlLcMMxHLiVH0lrAFYqDhy/A/NoabX4fvuIrdLs5TWbFeOtRukC3q8SpT
1ge4laLUNEEkjd4wtYNSxfM3D4kIWjaXkGpMV1Mg9YeU0X/5rhoHmnizOO0bwLDMZX7f+2G8UOkz
n1iWDkMpzlRg/Yu25hPj2VAcKEUqqzLtl9OKFvq2sL8f9j2Ql6CL0wkqYkiTFZ4jXEMYi8a0F40B
xlG6+9aLWzPn1qW8klFZmuYLUucFJlYxjubzgXP4gPT1p3SwFH5LZEspwtRNC+j3DgybWMLOX4aY
yqnYhawqlNkRBax6T/bIre57sTjjAwYPRvneOK/TXLuA3+0kqSIV4+Z2SqTV7UrD84imGpiKVmZw
/diIXJ64yXMIrl8CO853FHk2tDo6QuqqZ6L4BNHqMYRzBC3t65wZmiIqDWQQCOJtJPRJO6c2THQq
oNLAkoMwbHuSuEsBKlSKzOIC9gKV4gAOSIoXn1LI5ZvfKlBxkwTE1C4bN84x1FgZ6ouYw6Iyb+Et
8e9leP2C8pj3CQ+ck/JkEaZc77ivofdJSwlJqK85CD6m5erZal2qyfw92xxBBZ2pynrFGa35B/45
Lbdyjg3+vpvpM+tOZ/YJlR/QcYtRFwc2oXp7msaMpL04szcFmMB/06bXR8OSR/HmFmxYFRNGoE6p
KhscXBZY1zwuuBJOFlEWQmMhU7QhlJnzsv7HhVDZcQL2z+UAJZth6ACMb8uPS8AbTx9aSipXsqtR
8M55/m5zaEPm6yAWG5ooR5cAj3mhUtPrF5EjowBckN228d1xFE8a9NVgagYvoEQGGZQ06XSxiFi4
sHi2k2gLOjZ9qhpc8ZiHOQROjt5KXjk7B9vbBDxIJLRwtIZNNVDrWrzoBVg9utD8oiATfIGneBJ6
g30J/zmN7HNXmwWZx/b/FhxJUPKg1AA92vg1wcrFRNGULnUaaU7hN0JUbAzsT6wxHtFh5pnYdeX7
06OpZM4ojcIVMw4Av2qdTxscIqHWZBVgPHzIK/75tbai5H8DKvgeZcKBpnjabwCet67+vZcFiIPz
2F+Aw3gsWbNd1F8ey9xtUBuFbq7oAo2fSBv48HTH/1PFb/0szBd5XxftIaINtxG+n5Fdnx5kYaB8
GBf+oa+d8odGJgQmBdTgG4cMD6O8Er2+jbAfOVjMIneJv1V6AI2AvMT+dsu9m/4CB8XPZX91DdE2
swfIE5tyc2xuCiCbs4QRWIwKX2HvKmuXm1ZDbAyJh+is/DxR0d04E82/FavPuYXlfrVQllKmchc/
CbuddrU8hh3ftoXJ/4bUCQFvdSaQ+HbEC1WbiaWvudjQrIL2LWLsf1nvj2+8bIhX1t6PcQjHnL82
pevLkyVaVoihVFhdP+UFvH2UkqVg9p50P5USHD3Rsf9mNtm4mPt9hJFGM1ZUbog5uNwHHdOEYmTC
sxp4UjKCm9DJa3d2RiwYBhdGSkKuxrkZeAapUvubtyVRppTLecKYLqoSDtbTT0BjLWJe7dAZXg/k
YSPPsGPxn7isy5R1+SAf4Dbph7YNP2jTOtFkY2sOux3Ox5m+2L9tIvXvSTvBlxNs42PBhbWm5n3E
mWgZdMVvFjzIleVROWPRQ2KULFF8HRZpy9XO/ox5A6QaZHzqiUIUl6RieRu+H0kfOGWFfW5wQNeV
Elu28wUh2en7T5tKUUQlSd5ZQO0SvHtfnN0Y68smzGgkT10+iGESy8HLpyDWeLhNzXXCxcsIe2nK
hEO6gUOhsIbCNKSisKR4lQSvIk4WD1HBIcahKiIrU//U8W0M/4hgHjNWtIvn6g9o2pRhG1grWnnq
s0IX1w7QitWlF6vIVnpZ44o+9ZiNt/m5Sl6n9F3qoEiri5TU2gOB+nHUkDzrQFKNLmWKdNl1Pv63
J4MgSRbkr7jPXUK5B7Vikw4piEVqXOu5qO1Pe9HxEb5/xuyFxpzFf9kWlHL9vdD5jK+u60GhPcTf
veQF+BdxHyMBWvZkHig09ZtddCctsAqSDIsTaprCq5MzqvTqH4gc0wGgad8Xz3FU8RrBKlsfW7z4
41mLSlFSqiZYOkyHm9wUiYPRlSuTkPUck3EL0JeTVtofPxNwmyjooNVgobke89kFttyQC9/3x8QK
mTGFa1C5G4CYXqDzDwwXHb0C4EYcoHKPs5sHyuMyU0G+DZftHiyLh4kx+vs/A7763WZ2Z90E5qc4
PjjMsEHkXLxTwE4J9KUueCyKO0IoxnBITp8PT/0Sm9hMu8EOKSHTxv8JrPqSr7awke+ZCz+rw1Tn
9HkZSpI0s2QCgZCwG5yDS4sUk5/wXIMUL+OUhi/45K+521h1FkTlaCMTwn8cQ+an03JPkpy/po8d
iH0L1/yRHPSolxz5ECiItL/UcxgX/lIoj0kKB/6nVzIkNY4c4S+nLzBRQdEdJKYvXMiNFLm/9PGB
XAm5nuiUQLwfKEmvGhPS7heZe7g7Xcf+F8uJajKjzTX0Ar/1g2X1kqbkAlk4QWCDP+FeXN+TZNAL
O8Z7rOGjpHSKFG7XNMoFue+mjbEkCsTKodDCpZ3hpYGOS9qKv5nPJZVO9+sqfQaM81qZO9ntx74l
xjhFAea+v2Ux90JnTtKHyXOtbn9JImPickYN6u338vm4KvBr2f5fS+ViNj/MIhvgxjfpgEV64Xzc
NYSyuvTNtgVXJWRZ45JYwMv7qsPVZaL9MKd2xJUtBUmWG5cFR+fSxkroiiVMu4zblU7u1m8ynRYY
yiKlVLECglNMO2esLffkhY/I7EoJWWTFhE/eH0/S6TYo5lMrM1yOvn1RajTGg/FKgwZFD0iy3fEg
np79j75uukCrD+Hoc8SDaH/YWjhkcC2ebA/j8W8eR2TjXFeqfNPm98FnzwWmpGsw1yndTkoq57Rt
FQIqQfVQXSsYtz+MoawCFfaHcJ8kIdVEDpC4rPaHUkyjwM+Xt5k1uS1wwvmKrnGVPDySa7ZK2lLx
ZBbyZO1uS1qRcaz0KFGvIdrRO+2hXR95Squ66xh9qYzu9uUE7S0VTPnss5fO9gUv7qLPWOVUSIjn
4WaOXHKcryf8CkY3td+U7pFfOfleYwC5LQB7ZsuM5SpS1OMpxI3vaeXk3eTkVM5I842xBZTSn64R
OpxRXpv3TyeBA5nwRJx8ntNrN3XX/TB+ECfC6gWr9L8L9wAZuP5r3uK4X2pO1axeaCboD4RLDgLy
Jhk3zangW/3oA11Vg/jS794E8UJZ6YVFNfe/tFo8jjsVdyUfE/hM9CZMMjBM2Oj+yGCBiZmXhiaJ
AuARCxKazgNzrIjb+omM7ir15ImCMVEzpbMK4yYvZIR4tHV074IeQ/S5yPfULtN2yDmgGFKfi3Ch
uRmzDHf6D1HkUHSf3dbVr5T+7JI3aEADHgynvaCUWBaXtezm2Y9ZBd3MuWbqPeaKz2dnfC9NX3Ko
ikl2BpGix0e1LTUvpIHrBlLgkKwtTplY0IFz4dnMO8Nyi+njIuzLvFzpm4IArYB+xf71T+B3ySVR
EkLiIePfxLV9ASig/9l/BSTP27ymklIC6gP+dfdMyOH1LBLAvouwX3az05MNl0yZe/7VUyLnXQtM
7Lgp8E9u5X7CzXaLoXpagr705NolhZC0BWUeCZx3zm/dse6WglhiIe6eiPfovejJQiTfGm2drZqo
aUHS4fvaecMEZ+BkEuKfr05DQ3zye2bwgp7wUrEOo4xsp/wsxY3l4dPLvpZpzWchmKyFsKDQw59D
Xb3PoYrRg9+4J88dm6xs0fY0lDUISE40LTAazPsW8bvzCShIurGLvEzRD3U2dVyWeXuAvyK5V4Ur
t8/CArg0VKPed2EDvA58hzdCq6GUArxMpEpb+Yu+xs5hF0Lv2A4FwlyzgmOJL2fNYubeUk25GDdc
GO5FBec/Yc7xX+14eO+CJHjE3ScIFdHVjvCSLM4Xr7d+U4GnmYBMwMutjxHoCmU4QhTfUWOOC5mk
uv9jyf7enhhKxaqQcAfWRlUjeZUBEtvzW1PSFvp2Gkjz+jMN01urGmtC2Vp4DaS+KMEIGUikBx4c
rfrjt92LVpOQYJVrp98R8whwIv+Ibor2TDlve9884dzk6shIBIFySB0u7xwg2hz5ZQMLseWd2cQL
z3WwZIZiX/4kHDhibh+IMjC0vL8f7U3UzJwqxWgA2zEWhmWe0VYHt9hdiqvy+qsgrEHRSxkxKFmx
PuXZRgZRILeS9JnnJht7F0umiVTZ7J/kyKGXZ5De3UCg1PeP3oOCWLaRzTkA/LD7hMtqPn33c0J3
NauGJ1xL4VhJEEmlvgChqc3POR9/Cc5GdrdZNHZEnQPT3urOaor/ui0KNzCCFmyG8zfkGam6xiq3
3y9NqpJjkMdDzGmOqG/qApItugTIPuczuMQIsFTSd8bQ+lSPiwkHyN1J4zNbpPCX8jlqyusIL+iH
fCWuyafLjG7yHyUeJ5yuBR4klrf2kMTiCUrs+xlunTuGo3u5/Y5DG1RvOe8frtfBl1oGAC680yTI
CIe/Ug+T3KLYavUaMq/MmB9nVjWESc12ys+iVM8DMC1Qnl4ElbbuuM9X6bifKfGVRyAR4a9JgUEC
0dQfbkr9DfUdqgs0QQSSQzxy9dPoXHZtM37hisbm5A8WQ6p58yycvLRgWINX2RvoOnoksXaBr97+
40O15Bd/Wbv9RCe9p/5UYq0hfLldf2Z+0tGIuI5QyC1CImb0mdgKV0HAsdM8rQY20tTC5OhbbBb6
tk6HHmunjVAatE878BS7HsBh4L7/ZVKmyETTjsaenbnsdgq7Tsn3iYdEvJp+JkcJogoiP+IU1jyq
JfFT8GFHEJrBgdy86q6UTM5IlkxR/fTL5Z1pmZ7RTAkhMVbVKuZ4DTzlky0gPjR5YAFYFSAGDowH
9KyB+gUL9ye5mwzN3bYhf1mXiKnFjy+FU6gn/AYZ4ujnxESln3EZdX7T4AH4RwYm/9U/MKDMSLbt
NbCY+2kTth3PQ4eSe3l1mcm3QNSzKi15sSvamHTJN8wXCqQvKbx6n3eHBk0h+PuuHh21J+TaQB4q
Uf8fX/YuGmzZ8XRr40VtiztPl8+47ZCg/P+2HFHF5ShxgwwiTL7fHMfiZkU4bfOzDnude3b53oat
betvqCYiXJ6vEGQROGqbR8dFkvVIXQqnEIBSnQVjfZUjn6aNtcj+FQxy8OBXY+OPX8454xyddlgc
k7G1vasG1UPX1VRnTPOQNFSGb1n+uN8MAQBlM354eKENgT0yPgJBop6mclhmFhCCPE/GExxFhQCp
O1ubrhQUExbP5Nnj59ipqee0JIe9mKcS699CTakDcYBjxQQdsHZM8O4eXZNHP82wc+AnOp335WHO
Xa2jSNxLEnRZzJyxK5B6SBwspAfpTp/kK3q/ezwzkYXtHMA7B5NsecIBqyDW4fc3QWKbQQQ0tQuK
+cRURwARlBxR/xotrzEGXuLTOI+j6U3/17c0I9HIURlhOiOUFdNYuZe2Tnvn/i9u9oaBepwsqYp5
i4Vu9Qmlqp59YYHxAWzyzYr8cyo6GM62WMVepOJWlXTGkhzIO3G1KcfPzbPI2WpmxIXUUFnhT6FO
Pa3m4HrXfk9J0T3cFmfcXA4WvHwF1ilk/Ibw6L3Gh5NZqCQPN19ICvtubvWEgNX1xbYet06w+5Rt
5XUj7LVDL63CBTx3xi0kJOnN8Nk8Of82ISmMn7c+SO6LAggDioxACQwVEqr8g9ibVjnErqGCKVXI
xNWauItMmm/zWa+Jo2eMQ0l14oi0ITOVuD9bNBubr7Ej7VfGfuh8yjTNlLFnPvapoONU4OJzTc6j
EbJ7vc6mj9Z6Ttj3EI7ZG1ep9IpVeZvMpCkesdWnuMw8bWKj2dH7E8Flu49D6fSLidsKLJVsZka1
+CwsldzsxpbWLyMlHyC8RlA+yl1k695X5eLTh1r0uTPlYw1vQFNx1sD2GZBNt9STSf6MpaPem87y
G35wttcWa0kpDSYd0Uwt+1eyXFm0VVmXYed1ncKFrVWpZC64U1njjzbqQMaLfe/OlIKcon1s4Jbc
m6qkNPijjPohqDpUvsgz4SPoRzbb7V1swk8nFll8vE8/ltLYni+N+0ShZ4vQ3Z/ADzB9FkewcS/B
D+VY9Qut0dW9OpVLygQNhuRKPrBlG/f4R+igWXRwkM0cRInGEEHLKRJVHvk8EFXlCYt6cokBU28l
khufDrnKS4tZYFN9Cyhcix/LvWYCFFqSx4givQjuC7So9V25GzgyYD6P67vi56+d3mZE9P/vb7d8
hTofcozRWWWSrVJbGG5jTCj6eQN+tQZ3rkjLiRjpqGMp98/ATHe0aAuFV5oU4Lz22qdeHGOzv1zQ
HKT2ntMNKkkCAmIEI5+pMffZldTeoqAm7Ft4MT6D2jacL55wMuBcJRuFJ+lYQQFQAP6k8NqvWHgH
ZA6KspWS1Qg995Xe93FBpHO8M9T95ZqdQ5KGjEpXKp5N/ucchBcCFAOHYwbeFWhUksPPcRrRJdu5
TKj2+avwxx/1KaaJ8WX0oZEsw01/zmdQyVcIpzkMgBcOcvBQFDLi1Bv196RrFso2IJTzgcJZEDqg
0iVIi7MRHaGsJo1EJsP3c8n/KuMyTjRpplpWXNM/SAPdrkHRS9cSBGVuKi74FQPPJdY+WfuxcstI
O5OyO5MCswtKkRQ5gQdSiOCPklhVcy5VBa4PFwJ2mrnM3buKD+vjIwkhlsl/J0BJb1q9vaBBECpb
rp4p1Q+gx/9d1fVLk3E0bF562O6T2fImb5jRQlMY7xzBQ9QPhWuUT0U7N5qX/l/Ing9JMU2MQ5F6
Xs2oaxy+/5UqHzik9v7lffzC1RPdEO5fPmOeTlSituQ5TPqVzAaSlcRwfjOPArH5PZAquvPKokXI
WKP2XYHypXltvC50YxPoBy+/Ih1RNWdm4i5RMYNpOmAjCkVlaO9BxAjQYCXuwOXltemB+1ezLQx7
x6y5AFi9BUYpONK8YkFoyucK3ZJVIESlUILgx1138DlcC6EPQYeo61y/YDJ+cLf09u0ENSZMCst6
hh36VfsSWoP2itMPPpEx0PUqjILqH874rAxfr2jb23r7SwYwMGhgNAgcH6JSfczZaWZyhB3vTtGB
9BjPMjJ4m5edWddkZSdc8wCS/gnv+1bKAix7JYCei5HhkHvsUkAdLXN16NCqibKLU1x3QoR5Nwk0
r3yXLPuncAPTZWf9thIsPQbSx9yPfAOsZixFzfu7Mfa01skpl0BrkW4avsavxPLG+/IFUa4fFIDF
7IhUXaPQh6H9ghyH+m13nkAd5sWFXTtFoEjc6pzGdix5fr29tkWXz9/NkPyEhMDXtniFZe9Jh3Hj
5HAP43u4BHZ7G3vzdbXsF43HbqB7dpKSbz8TWvoN6vFRznKi+HgYxb7aboQqgedkPL77vACPfo43
scfXBTYjMpXh/UbYuQ6BjP54SwoHxXXU1xhVW1iy/TxbezU6S/CtASgbc9Rh0VF3ewDlx/5FQ3g8
jxucWycFFjsRvrnkWxIp04+k37AmRsI58ERZB0nMsnA3O5wQEmHOxmHfaIgM9j7jPkjNSiPeFGkP
0pb74U3iZ/ta/Sn+3H1Fl3lij+Nxg+DYHex4mfkcWk94A/bQ0z+CY3V7A/sLu/FmvEnegTUXIs6K
ww3QaOD3m4teTMKTW/iv+qbrQEMTU8U/NgUe6/Z2uz69DhqhMYnb1nrQEnvvvto3Zhpl6GCFYJVz
4pQxX3Opq4yP26YDjX0LMUhSe3q9O6Bddl0GrV9OzqfJY3caEIvGsdqjF/CnR0fdPB+U23kde0Fk
08xJkYsAqVCrIg4KS4FxWUoppfLH9NdMKivpLcFuQeffFkSgNvKMdjvB16ILCXd8afPhlv0d1wJm
EC70qJOHV9ZJPdyfNfVWFA00EgSamge4L7hSgSXzltUIN/BA2VeJSGhET5dWGmpBkFjlDCbn3IZD
A8YbvA/1SKnIp3O/6SPxDm/NrKPbl6tRTET6Tyq1TysK22XfJ+t2ivVxVellLJn/p3UHJ1iy3en9
rAzNCsX//Lsl5ja4DAlPouLisArtlQxVQkLZ+wB+c8MviwpQhfth7Sh6EVFwIsTlvvU+W/h+AlNv
qSAxHGYg104SAR4ZWQs3vueuGUdGiPnarPg6famR6oQiWlEQXMj3f7l+UZh1k53Vl11RG9BHydMa
SdVxAtkbTn/iDWShl7hPJz9wj+iXJO8pSh9Ek5RicwWSP4GQ3RSVZ3TbxXXmvUnVoWd8+ls56Di7
moR2DiTmpySFCfuy0iruKiVQ3pPzh+1QyFhaIXruBSNuvSrB+wQJk8SuoEgKd+oD7dWonU3cuPPi
LoQlOpOZBErBQ9xUoUt1g8+LCHjyFEfXeDrKOfDE1ISl+om9JB6lINp5/YZWS7NYOC8TvMHmi2yu
JdZbgjXcJ8QKzHv0TCp5Da7T9fl2j/FAejygZhAgYJgFZ2mm8b/RIRPA6bjNml0RlZGx2608OCOb
lwisBxc50+5XhbpdHHctj3nAU8TI3Hcvsp89YbkQtrqlDgh3wftESVSQ05UbGK9b1gL7u/yBxQXm
WPBVHFVuxmMe8cF4un13G/ALBUtqcFCvvaUv4h53cRZc1ysSk3brzf1jr4B+dsU6cGbSrePLIBEk
W2c7LygbjBM7rCSW/MkbT5UWCPhowYqMK2ApXF/QccorJ9uBjOMUTds6EmRrl82X+iI4sU8ifI+2
jfwRIqCKi2NyT9UXX/9g2HEvdUgd48CKAPUcP35WYqZw4lmghUA4BCLBMIKPh1wwuqYTAt5TUgDV
C4abDfbkQOQbTpkt8LDy9Oto30tVSoGm/TZ0fW8DDHk3YgsmSwxxmW8f/ZnLFLPvK6guZAOMVt3X
mzmGr84C3yqHXdKIFZ0pRRZ4Zp5e3LOwVDSrcp0bPdF8KV/ndNoFmhncvvsxCBd/QrssPYr7DyPP
COXWOcidCK+LBe9alNdTNlosw3Hwec/vJLb/P0Yt9qtWXfiRGQ/Thiw6Jmrk3BhsnTL3c58AYree
83CyClTGxdWVuZf0u0reX7hphv2BB+tuuNYCuzUAfl4LzWAouLAfjPY7hMit3a12Zz97oc//i3Au
GnMffXkPyJRenb73lgqPw9uLvBgzo7LzgBrqv2mQiGdSBoh63HjrcWSXBFtyRjQNTaLq3A2qQ0up
lFztsS4ILW76dzZsqd+hAEs68RBxfMpTApvxl17SzuVFYoQ9B2IKiTGldysaRLR1wzoIXIzmQ2v2
1Y9XlVE7Wv++lMDHbmIrYnqMDELp0A3TbYPfZbTS8ReWvZuibAFOD9f3QqINGD3bpntejr3Dlkp1
I3mLo6oYJbtefckJ3vk+hpR+E10V8VWh5nz1R89q+Gffb8n8PAanfScBAr84CtFxz9HCGB8V/qPC
jIbnR8EoAnYvFdv4s3KzpBx6A4d8FDsWMiS5MaVP7XgRORfWhWj0vODD6oHWxXSMBr4/vnJ3f4xR
38UkSNXp9dkZ4udItFM4SEhITGz1ah9w2t3Yq540drsbOqWSsf8sUaQXSs7/vdEFRsS/6G0uHFN6
yFs1IE08csUb3Y27iGbGasWW3hEWGciTYDaLrvKuU3riyBhyOolF59zp3b2STO5TfCQ80jkcxmuj
QBiwbDk1waXJyomMBStSrwJBrz465pUY5/XD1BRFrd+pMJYLicGPkqS7Qo4MyLFlgko4oRP2jdnl
ioRO/TW91p0wi0xhgEUKuFds+EhxL9AMd28NFO3fZjoAvyFJEANwz81ezzkU7cSILadKmDXp7I3/
TRiwnDFc8I6ojRYxEkEjd0Lhbm9ni2BoDHhfAtRrFZLamD1ThQQOCEIn2whQ1T5XQ3U/t5UQvFn2
t1DyjyYXIpTUW/q6aKEWy7K95SUTTlGfmTNY9ptyz7/mEDVLPJr+iauNKj/tMzTnFiznqEBh2btt
zunrxhd7MQWtjTujogDqYBIQinUdR0jWVluc45B04n5Fg7u9b0oTIzdflsHdPjW3dMysIIjDfYEs
MRXUilA11uZwz8/KFBq4u12XW93KLGd0VrJEMMpy1Qn/N4aV+Vc+EM3sh7mS1jeOcTkR0rtSXxrt
RH9lPQhNmWi0R4pSmYN8cfPO2qDDspM5nfwLdQaE8p0QjJltlj7JHYeb2w7+m1ialj/0SFs6uJgK
QHVwszWF0gXr3Qz68BLrlL8oQKwz4X0tk5RgmsdB5gSj7sVbWgNs0uTTfG8sXz/nRtCcHcfYerXF
qnqaEQd/qkXa135gZT/yN1bTOscxoQUFKRG4ceRmTEwmmb2wlo2WmSrBHIF6lwIIoaLdwc8mBxFM
bMk6SSNi33fkyT0jgpW+TG8YaCL6GuoT/P8a9/q4waDngOdAi55IMkz+4yV0mMkVYE+PfH3fKTX3
fM5DOIHYMjUBqgp1MZ2IP7iHJyKQ0a8E9hU+ABzBEc8afAEEIyC00a3VTGXsP7DpfW8e7wObo63S
x0gJFt3JtGqertMZQAv/sNuVhpZ3ZoixSlkxPYUy8mP/zBoWaQL8j75jDKLcM+FRR2VqkP7LW6JN
YWtR6Qt3kMXyiglV1/X6thqZldGY1DtI7qAANNCqpKrcuRp76m7ekKPSyIW9axMalez6T8TUHotr
nS/EhluwwrL2bAJQa8xWMNn6ze6lmWL2QSS9y+t0WJaC6zlMn81xCwn0TnET66nSrni2M5nL6Rgx
/DcmPW210CjbVwjUWDWwhAWzqkCvUT//2xnBpDNh6UzlWTqjLnwT+B43aS1vSh74hWpXe3saITsL
Yq1WxGGM/Xgjkz739nVZM3EuNk6N3EOtf7MEyww4bY46n/5A6RGWgbvHXLc6HiLRQYIctdlcpJ+n
Wh96Qq6pZnWBpRYFTGwuK1IOFKCZI4M4uwaNWpW2t+eWwK3DcGZ+OBuOb3o6UvRrJZDNGuAJq2yt
13DCX/5UXPEtA2Ax7Fb0OVVtGLcckFMiYgsaZfWlNwOgpBU605j37k44gFOhqOVsuVVylAIiIK46
EUDEzbdnyW7rQag2mogziVTFF34KSuKwBs7xjjXjj/hiOft7lGLrZaTL3KYCN47JO75zL3zurKYD
BceTmn8SdX3dh0OaTxp+MJ/jyDZ0bkh4z3WLhEkLHqxyANS5yfPdt9qxqWnsYn3EKWvbuvDOBXAK
P9W6KN7M0pPCWecvUbnyZqKxq17ClUYCdYvTNtfJVzS5VpMTf10Oert/eez+JjFw+Di5CpR7CQXn
KvA8teoZuuLBUWLP+NsUcKeG4VXhDOTQABD2SL4ZzRnWa52rnQVz3oHgLaG1yZgfoad7EJM+6cvF
ONKVk/QLIZtaYdhx4bW3xoPrrX+bXToiE/LmgvOJphCIp1srwx08m7ZNp/b8TknIhzHwIxF6/Qju
Xlq/i43jlx7Jt6PqbjY9F5mswDV/ohW3c2nA858SV+nVVLst0f+afwNd+MQn+jVbJvZz5IPglyaY
Rw+SH+slr/6gMBc1QNoriezYlviJ2uA1XBH1QVk4+KX3fGWfhSXIlrCIECs9Qz8dEwMBwbwHrXWO
RTC0dim2dTKm+SL0bJBC8rDefZHpe8uu7+eFdlDFQG8vUA/xLKvOs++UpqH179sG/GV22iQwCiLB
gcoTivi3FgPVfVxSyIEFktxRQ9iwd02vTFM8a2WU3mh6z5UxPThn4VZrSCRjP+OkV1fmkafH0s+h
QOGfCZ270cmI1bDMNf3+jg79z0iyNGP7cV5+3eLqov+ubbZnu19/7+YfdEMRMJdNmN2wplX+KQ5x
iQxEpPGGWS+P8ahCPd4yBaXyu9UXQ/AUXLoKrqIyIBTf8ijT84XRSEb7/H3HXeyFvspIsg9qj4P7
ojWAzajXGPJ/1JGAq+a6A/oFpAbI+aHYRhqsnVFFxNHgEz1R0FDmQnoNrHHhDPuCiI2H/GHOP918
mlFoKA8HrQoh1Bx+H6xxD8c/Bdu+fJ6DIIJK+B6uKc3zg0DIHVYFeRCRmCMiZTgIFjDmCBoPzTF9
tMrXrAykabD7Pznsf5PqBtbtK5tc67UkgTY6RrmWOtAiJQnzY2pDz6pRquCWptBEMB68Ddig8K6k
ZphMNsVd4g2nITEszr15bms8WlQD/C10O0DgapKhDl9lpGOLlig7rx008wbz04SRwFKeiQuiegz+
n80TQbUT3T4MW7F/kwPrX7UbzspBl6Ywab3Xnzb4Gjrk8X1hjXt2TXEsCcKGGMMcbZoNYoF3lg+J
Zy45/KPZMQJ4vjfpJ/zX7KBFkRpcoetVeRhAlx9FWViQhXDXXxLAOyKaRRc3eRxRxoQNg5vkl0uB
/agok8S65ddV62okh+NA0LvUoynixLcTNiv6Rfg+Z8f4TrHw5UiCyKQ/YtJphXmS0FfDyel1IY9i
Y9w8EgRNJZhJsaJLVxQMyqNx8uHd/7DkKiqHCHkkoCR8AUcYhMHrnpivoA/hvvQ+N1wrmpBbH88z
XIR/OUTYm7JQTYo5w335oeLNKnM/EpOa/GdT8Z6I7l5olMCcmcm/b8YpjrJVNArc2g3DuM+aHXRI
EBx+NPpdXvS9SHdMsnUpgqtsrnCCPu+liF84mVngNEGqQ8YKz8FzSnDbCWzPbTc33Dm36lAzdlZk
PVZwUmYvcjnPbEcOj6z2yxSqRvz7wQhoJxbnt4F+QA5Cv7KcMoECb2ieDD3VBM8qVcyTf56lTnAe
SPDC5QmEyleoJNMj4nV88NBwNADeFr8Nlso6uQnGm8kRrYtrpF3q5AipwnEYYrKkUwtArsT2IsnH
OgY4UCOmnQNXQwgCIfkixxGM4W8SpP7/V+LMy2QBwUkYzLatnZlW1WRBGr1v8Zk92C112CqjDRBA
iaDJRKWQKxbGDF4VbOpgSCZZZ5kAK3geMUb3wUGNasl4LGaHqRw/sqyoERk6AP/gl4k/ECeTCbkl
4B4Gnesq0bgaslo4VqIiAq9dITkifBw1snvq1DOwEOu+O9qo85Ng6Rqup3Q/t72xaxJ1LwmBrtcu
/3ocw1CCJ1+ChkLTsQ8+tYNwmyIpjKVvTUP8IYKY0Bw/s9U8Z01HLGnODT7PUgOWI0MDb5w+5Kjo
DMRfiDKaxDG3KdYJHBdrTG4lnshywan6cXGHLErLlBDQbHQfMrOLyy9U54a1TLd+dVxIlSxGElPZ
SgjaiNaQ4eOP1eEGqYwZ2rWJl0+sLgLlO1AdVfba5r2DOZQC/dluGIYhxYEinrxZSp/wJyFKQD59
BlgqaUC5QaEfNXxwyd4EZ22bMofXk5ChI9eZ7ePrzRCUEu2I2QoT5Sr0glllG05fCQ7BP5wKbqaH
RyvVWMdPB9EBl8v9dV6UWwomcwzUOqviiTbRJn9/9BfWLeuRT0fwm2292nr8HBaOBzpIyoCgMyEB
sgzsdzGM/Q6ZZCMCs1aP+IvWxqVQ3m5AIQqt5JtM/eLYD3tyZ1RrrHg1IPJKAR4DrqgSFqX5L9cB
qUT1W5vGqZL5H0puuJnJ+yA43pu+vpe434yQJlA1USNaDZ+BcDMYIWwhYO9QzhcX+o2dHKlKYATi
m+c/mbhALJDlwhnTagYOyD+mWdcWjPcqJMVLDZp5pDGuRhBKLLloZ15+Xzj8xRXhDGh7bOqcRGso
dsQybGAeJIwRPFeUdxJyynd9QnO4DFROdtY6PwrcsAave84P//YeLhvZfkiaSOLZiGAYyAQ8/+TV
fhr7ZfroJwoFQuhgdR1hCgETgKZc7uPYm9Bh6oFtQTeJRKjAbzKmvoP9Hh+kXfUJ0FOCkPr4Bj/l
JjWFYvhl///xFf08jEqoZskjUweJTNf2T6GKwkuZyYmB9wtXsTdcZQoDfLQJXzr+tWlXnFXjtnHg
+icgL/0yfo8fKe3xnkRIc2vWJgBRcmatmZvzwYjiLAzr2adHF5LWCvtzvw9W635Gs+yQbLHUrBxu
y3GZdj3qxE/5td0wAHEY1vRUd6dB5YOBzhEJTWyfQaLNgIBgtpFzGe6dF5TglhrR7HDkhJo+rba7
yXBEr6UQK1W4rvrd95YyBi4pycLSEoX2JhxelZjwiM+ncCqpAncvqnajVBtfKXIEvRC6q3S/6I1o
pVMxSu5bfQfkcKjz5Jyzva4uXgSWLGuXBZy7jzV4CMNm4agt5mXL4QcDqJbP8fpDJD+1iz06y1CB
q9VTu9ewCV9fHEBzBX+ZcYp6juMdZHJQZY5oN8NcRkNEnB01lYAj2FL0VinzYQjeDQTEJRd0Wlu/
Y6EJyOHY8KdbMnb5+pWRYqF05udI4pLFX8wvGgxqydM+SZXpkj6l+lQKS/Is70Bb8/iR4ukJqEws
dfJ+QDHNaBQ2fb3MexdB8ovXSxMOc9gvrLLFW7brUS/Ua5u4GhPDnNs4lBUDl0IijWFCw2xjgn6M
UQsk3YS996ZOZ44AqIRHMavXMlH00V6XxzqMCBXMdGBqvk4oGa7fRuBanh8r4+cNTAQg9g1kfM9/
/ZLxVdvUXAp1scNO9LaY2CIHy708zjItnW68v4P9NwZ6LDSiyN4LrQCvonVqSpc8tpicKfKYeuPb
Lka2pbVcEPHL57IHb/1Fe8V7x8L8DaS6WyB4trpbkqtPDLe1Y60jXyBfD21uxSbUiF6YKuqNiChT
TslmcYIiJYQ+netd4LKhROfCurnvS5Cj/vHSuKK/PifjRmhJec1+1RuZBLY6GG+A9+g5Vzt34L4o
mUyVvoknJBtSRKuoNby092vsIwu6JgIVoz4E7vnv4aqFPEQBIwsQtmDmlKiYWqZAIlDJR5yhkCfg
SZdjaB1DJRCFHUalxY/KzThl/PskD6SRhy49Yr0oJUaB9GJokzYadvj3FJG6jGfXbH2HSJfBm0iO
mzv7wZlt9iXyxLiDqE/Sr1rNbPfdUZeqOKVamPo5Iz88WlMFrAH5bfMCYfi3GcUS2+Rzh7ls4slO
ORo8GokfFia3RWDBPtgBIvmQ7XMywxOgKtDrh74sPLrfZEOPUkHoYWNNxlHVsiRLJU8ts1ffadbV
l4Gbump9pRHNAblr8JDXY9GtVzhT2/FsSHyg+E1NlVtt+2ouJGBmCf4g9VmV0OSE//1Acseyoh77
F+vzMKTN6zPsTBTE7A8gnGPYccHF8v91XBMtcDpAo/wBe9r6CgwHvXzVMI7v/U+E/O92+fui+2eN
b2Xiya5m69eWNctu2kQivou6b2kESspFpkSUaZikfHiOudFkbyrNrYNkqecYryqKrzj0UNY/0B7s
tWzCFuM8cOLc4P+NKv0LrZh325se7P/IaiuyVjsuLnu/y7yXuRqxrBWLcWTOTOLmskEQPxENzxih
C+G0hV7vMshnz4bElg77dAl7wPOZ9o+zzzggsHuAfGibEeRbVva6qh3MGxu0kcVOC2z+Ab1KPxWv
KzanV40s3s6ptjJ6t3W2Hp0wuWyJ2UC2/sTNmhi8Lf0Vg1nQA3CX0m0bta+BzUO2sniaU6tnSFKG
k+g7URuXxG9PAS7lOZUfuvc8SwdthcMuI+34wcURKDBA0JmP11lm54EthzOib3EJ6pBtync0wR5t
fqFT2Xm1PW9U7KVfNBmJkm1vzbsu+nSVKYiRopzBll4IWxZM1Ec2snutFxTbpfGSHxTdUW3x+AKT
q2Uf7ggfNdLbpY6CoRj36xq/EUb7nt6DOTdULkN00jef0HSlY1r40pdiAqN120vOzorXp55+BT8d
du2ySV1m7dq2sJ1vlzRPyrcWGaW1VpcMYDiYBYQbhCOobzBX6cs1aEejoNHrOQ4I1l5OqUL04sST
9ABY5FBxtKbKPGz4LD39mlM64EaeWD48cuhS2KRssCEybEj3ur3RKV2uDSnwTkhMBvLw6ofKAxTs
n7FTenBt9xLWvOI/EQzMwhph2cjrzSOKM/mvXVR5ax3bLl0aQWFx62Lhxhk9A9BADSJpt8b1xJrH
sh/hqGqqIgIsQ4nMCBViMMtt6y8k+WogxgQS5pP0tp5ABE2/An7EebvoAmsblnTqBaN/Hgeothtx
3sNHokeGVYeUh3G2DWQEiC42VCX3gjXRx/tTQlPtjglLHqNTyY3IniSb6n1mLS0UFKux9itf4oQu
sv7oelFT2V0zoNc9Ss+BrTovf3VxOMdDUD+uRxCu2whhPwvQMYabfyal1EfUVVB+H5mb15HiC2JG
gzGbWDJ2ovcY+qZFZM/advC6mAtLZ0Ap/0UtvQkQHGNov6mRSjZj/DnNAqgvMQdc3SWi5TDoLxTO
ahWQI7vDzwkkhAqfH3y51DvatEIWODrj6qXRArSoFw3/vgUUGiA82dHi8Yq5cuQPFjGcsFhoPmPs
+lBwhSqRGvEL+xyPxy9Dwc0Xi1MAUkXykyszf1gfS7JrFtaklZjEZriz6MK/i71yMRdNmnzrdQlQ
TcsGbiied6gooulkVCyknzQO6B0hzolOfBEA/cMy0SAW/DnOEX48T4IGksK+5lgnFU4QOdo4UasT
ywPmaOVo2T5KT73HVacuZAPkSGpu1/R9tc8XrRBKhe8wHY/6G2A2Q40HXY47vTPgoB39ERLrNw+z
aYm0IksxcqKqIwkPOAMXtxJTbSCg8kdKahsD/f/5DxPM0izc/OXlpCFMFuNP3288hjmRAX6DfYyN
yohS0ADuyMD/rqq1zvWxA+36T3nPrY/qtMflutVhaaZqcRKjaczU3TIQJKJO9dfUfyr0WBeWkIrQ
Z86pwheNAM60wvKxD2m88rFwJn0FCMUTOpJ/gXmr7uwoW751D0QPcc/QYwqjjYHu/hlRsWOU+XSn
jTf+jopzuMrAmueu/X8rEnrc+0hOxumSfqFl5bYef13nKm+LRlX/rivwcimwMVcUcrznR8+nhq2l
6FBWGJSU5CCwcCygNOwKoI1CpS2xK5EGd3aEfVKtmkr8qzLNbfoznSq6bfvehBMeKf+7AcqhwZaD
Hhv+fmZe/oTFAerJseJCLNpMWjfBo720BhZFitxA0OZ3n952BSPMEVEy338wQF4i7Q1Z/TOw3AgR
rJasJIl4XOhIYbO8m7CCus01oNhCLPPwLjVrNUQ6+Lgu4ziPGS0ewYLFGuYgUatZT1R4a2K8q4JX
TtV27+kiCWyUiuIV7JgZvppDA6jryF0Gkm9NREoG7WxjRz56WpYKsy011GKGf0x1lEtAJP8vzgfN
5BnI/9KJWhjn2Lw2ENTLlOOVx4L/KU+ezftk44qvDU6K6dSxixL3yD1JMzF/bdKyppw8bYWSlQZ8
Ugt9lPAWKe+fgmEvsFkNqpW+Jmy0R7JdEtDCUMKQeWW/Wg2J+GmFBu0Huefzgk0dcj0kzxiyySc5
Sy3gR2QDjx6bU5u4QfcWgQ7Zo9ckF1W4JzaWAFaRlNSJCZHxwQkULMt6qXiKXEteF0guckWlejmw
2HlA4pElhDWy8xGrWyCZ8PVCkGHBuCCE3JUe2V2+D9rlleSD84rcYEHmDifnP3mmR8ZSOxyZrN2j
AJEwEbxOynIjtK5Kdk7b9zCs3tHVpSKt8e4ccSicXtdDyNXUwuvk3G3AnvwVjXI2tJzH0UGn2/FB
14sSxa7FiLf/JLSVrxeo3agGh5RgRBjj94Ywg7RtwoXsh2FFdPhKnLMxN1J6I0pjrUkamZIKvQZ1
oS4HTUYIeBV23cTsM5rrFAGywrBbLat1sU3pGSsExtFAKc8oMXlwkLsQyrryJpcY46/CdlsLRxmT
9Hlvan+OTEgU/zcPlaLohKfjOLxI9eDlu9SkQ2sQouJWsx5qqbZauJGkrNS51sQOvyIJb43TiPVq
D+jI4NLTIA0CZ8v9CpDw9yFI/YOCP+RKwAz4NLhPVtQZoknhM3/4HApHOMq2yYwHUjZq2x4wh59e
XR3/H4Idw+6s0z63qcSNbly6Tu03xxjynBMUyfSgStqiGnUklWHKMqbnauN2UU2KdYmSOe3Ysf6b
v1UzNln8LMsmYyiYG/21A2jjNWLgTFNkum4R13bE4nnzvuS5Z3qtYcZSgSJeCgZCUWCf8PI0CVcl
DkdAh3u8nHjvdmyBzyYJXOY/y3KNMVO6VF1BmExNDTBxjO+JzSsTyvlJozQvw08LL2BKDP8RIHq6
uDa+njXhhXSTEvmjpoT38QAp3t4u0/gqicTXXXBmEwLDplQZQbSdVC9/yC7NKIfTKvP0gh7UPhnp
d8XSoCxSm2srn/ZaVUvquazYl6Cla1lh5P9hahZcQWCYFoXwuah4+e6Nou+Hz3LBVCA0tWKsKhpW
tyy08J11p9O3Wis8GlXL6a5/TDCQzZwx10fudaarX+XFXbrWuAahoEL+oMTUxFe+gYvRje+JYPhb
yiuV5BPcudJoII7JqKOOY/aFMm6j/8WAHW7Xi6LYX8N1JJbI4+iLW94726+3j0c+MfgZmDcehKT4
Zk+yFZXRqvgO6Sl9c0ypa3gAPdi3dXl0jq26rwf8jDAeKNQ9wjQF+aqjG8mKbu9OsLdLSdJL60pq
9a8Fxxu4LT3NEfuR0se0HYbchHKFZmK0+Knbd0wWc3Bm6TaVHqxrVuZ63Ls6k0LWI1La+dQOvXMF
F7tl93cf/aRjOi7HBG/PhzVREu6BDSSRuveIHwljAG600OhpmI3szXHm8zyLsgqEdxJxTh41K1Pr
NctybqX9hQMm4NdxCMJBIDNNaUWbrWA2zMjGFDY1EzGT/2lBFPbjC9hGnN5ciSJqJlHZ1CPBOdMg
aqQU721pUm4C3QVKug1+VYlT+bjGKtgpokbXd3COCAqSTN1DUESwQfPoDeXjlq5/eYIxyOOysSra
+tO0Y0goZ7dLajtI3UqMqpHfiIj/MW6tydVHo9TJxwVTt4A+J7aQA2VuqN7nd5Xk11wTKkkJ2jnb
rWI5FBX3D3p5R7yOR6f4oS2AvGxADB4zP729V1q8mu9gmNCW3WCOG3JOzKFQKgi6OraFDFEzrMIK
V4EqHGeubnanQ9bQN0Ppay5qUeWUKYBFMgHkf/Wf4dhDbg/qiHi+PuCdfSoY81hcxOldyYqC8y1J
rQ5XnH2a2bjWv2ZL0x4q0yaKFigpYkALpZAK+a+cwl99156Coa2Fh1ipGABTcxdmcqC/7kIv/uf/
JZ4ggxQ0JwxOhfox9KpxqnCAHkOo8fdJ24xPrm1/6WbtB3CKFZY/TAYlLKlEKBUQlVfD1yAf/JcN
AV6aq4GTFKryXsTvXi74TjUgSLwAH14GHqAD/sk44W27xyT4ke7OT65OZtR1gijXID0WnWVAsIFf
sjeXXaj5g5pQUfZtkbyQ6Ad99Xpxm6ikTea5Fs1LPzxoLpK3d0sYS5pjgSi9hmEEzbNRTKVkqk9V
sh8HD5kTaBYJI43gP47Qo+XwnYO5d61jQfPZzoliE8e2OGBJsAcLieJiFM2cECuWdiC1kw/Pg2GS
fEtPtXQz5yCHmbQkUy8UImUL4WZHjhrEiDzOmrx29QjnkDkQHp3w2QdFdOmNzRVirA0tfQGSmRxk
XVcMMsnTDjQVHrvldxM4pbTrM4wazyjr+XTjB2AtXlBGh839TyAzjkqSPmHTvHMUj79SarZgY8ra
xAJ0C88c1cDPGITE6DDYcKjCuDW5F12AIunmpPS++Q1Knrvut2roOXTE7MG62pswVi78A0cbsCyl
YUBO6xDeXzjzKRnP7PcJ6Tsf0mLh4ZaAn3QwvIbq3AhaLFH1UHkxW/z1uZXqf9e0A0B/GdmL6flU
Z3NQ+KDHCWBdlcrKT5eNfxtaPWH+ITBy/t9xTRz2aKxgchewAeBycCrfzLBl35mU4QKbm80OsGt9
Zi5zhHvtNii9tsb2C7C3nbP2TWBbcHnk9VmQQDzMVwkqDxcnVHz5tEPjyPcLtFqc67zfkifnukSg
K6B50lFyzlrwfFQv+MisejN8lExNIpzRWJ5hw/P/VpNCR0djUdGdLwUT9Rn85lL2ZBFsrsEH7lap
4i4HDgtzICaltklmRK7sprUq6bFCPkxV9Ja0QKp1TQMLW9BMuKLI5dGxn3ym4/cGvxY0mLPvvRmX
BcgDfnp5uM8rFn/51S8XLCdhHIsv8m7EvDq6oDn1bFdrkx6omLUuJMdUzdYgj98dMHXsJezOI3+1
MmIHyEqVEYQoNilMq1j+GyTGTcV+5nWPUWUFqYBtE1Qalg/xTgzcVaBN7dVvNm+ZiTDeMXxoBL27
xUoSo6CjU55LR4h7gqZChmg9DBbIqrXFq+8NnE7zanE0UtV8Xs1l1diSKXrhCoYmdRz1sBsHO/3G
EJAuWZy0yph0QDxWrf6mAk7xtkscv6bYdPHQbvXSzN/oRB/JSYuAIUftCApzRB/a+eNOX9RSNvU7
jdrDsTdLHAeFDCMMXdfy2l27c0c8rJzjH7PT8Lcc8cpe0KQkgZToGKDAstGhIi40hT2rvlLTQ/o4
9Tg9mLq3/j3Sfi2D35+/hy3GOSyovDqdlLuVvwc9IokTCcGSR6kjQPCB8td+dND6Mzw/X8y1uaVv
0TAZkvb65FteN04HaheZRoNek9/HjMHndJN3SxFSLsIP+fmFMV2Tp7ljt1QtcVOmkE6cotdQnJTB
uHMeQG/zhvU2s3Xyrv4p7tyNRs0L+nVv3xxtYtLU5M0bs3jqZaCcz09UtkOx6W5mgT69FqIZvhMs
yZGww7TtEKumWF6zlzQRnSs3CkS3JBFtaVHEPmSxzqrQ7Jkh5JOO2PRqSIdj0zbMGuVYz4upFtk2
gVXHBYIp30hM8qbj+S7irCvCLatwQLznQkNNz1uZkuATlTkrnZL+xl3GP5lDI7+bidfQBIrtmyIH
2Ogm5PtwisXIO+KHfP5E3hcZe4sqPiCwlQ7D2P45WzlR0ars/EOAg83C/VcXHjeI1eG5MZKSbDi2
/+GNl4gphSlJ+HDqCVOhhXnL3JWfEqsl8ZJvLD2yFjOd8xT8SCcy7yGN7qyssSaFn1FikPwUkhiT
ofnlgHsO+L78Flnn7aYzOx3pq4nVo2PoBTN3mxLLzLxf6BGlS0J7OhndXAPHxSgvjMDqPlLgK28G
vYCsdICDlo/9LB7lqou591r/8G3+3vRFppH1TSyMhFx3sQaRzp8SSpnQup68iYbQSbkOD8KycIzl
kVj1fCNdgZcCxzr8kTpxQy3mpZCcV/8/EhGGM2F9tP+4QNxQb8DBi49ZJp0lsPD+7tQrJrFaemaA
RRSb7zFrN+ElW60NY1R5oO+aqgL/WDdEtLnBMiGpQpuKyKbjnUlLEE7YGRGn2pl+ypB37OiqEHDk
7N8XzF2J9eQUABoVj9I4QLQ+baxVMoDH6Un9BThngfH/MuoB63/O83nD/9XQuEG9NaOj8EjQOcu0
9kIoHrySmUyxY233WxFcI8IzLF7mPubbQjeLKh7xRWQ3rQ7S3Hu/hfrGsiRT1DrAppwugVqVhBSL
PyWsLTDYdgyd+Ny3/1L53AAC+pABG0H2QCzokSUwCbOXTE/C5QHkr9/CZBN8oK4ppuXJudDXfQQa
/Fx5MEXFsmYExJfxAMNGV3F5TTpHF1UkLHJsGflE6lAM3i0anFW7Zt21DCDyAbsDYGBfpUP91nc3
ifRQbihYkQX6QBCO9KfjAacvmE6UezKY2XOKdOUDirVaL7fuIE6FSnh2AqiodAUgzliN7mPlM2md
z/0RjiJFgsjg6cqnJftZKXysvninExlcpU8bO8ZiX/30+Ng2US6E+6JlgDvOvTR2qh3gxW4gjlVB
Oav3n7LIZ60ZoJQ7h+fW9eqzAe+9C0xbQb/WptxdhNi0Kh3H1uOy8v41YjujK4RjZ+Sh2siTEpef
OF0gtYgYmmqFyIGEvjkX+uxlX+BKxXMCT5K3QWaTEJWusy5eFCciJBC9KG7bB+0Ie1WoU9X/Y+D7
Jbg5al/yhN7c/oToL+Tl/ni1cxafKxFWeubuTjYaFaivQ4ZjAN4FSsWuFLxs+MtpIXGn+rAy0+qO
6HYLN5wJGye77AgAXGXuDsnTEu4temEX8zzSLIIMdIlUip5ZXJLGXGhaq4HNFpkh34SW609pGsqy
AeNFQVU7huiBzbkWZ12VRwctr6VlPLpqiZakCOlJxHxPeTJydN7BXkCST5OHtyr3C5Yu0aQoEzbs
/KJVkewsQFYKxvZChgUp9rkI5LxolHakFvnLqI8sT8Zi2gd3cngMK019sBFF6hphxVKwCC1gEB1Q
xq29AEtCITp355C8aYf+n0yqch2RiFy1l1cJ13rwQtypzLjyIXLAm6oBgruIeK3DLRAfUqtjMyln
Xp0PF5UzR5zK9CAb9yej7MJlMKcDyXXea4NwvsGYgrfcKtmbPVyd0BP821iMDbeFlZV5s9eZtnw2
KhfdHrFaJZC+oVNk9dB/HwA1m6cgYCoGunwDsksLkzxeNGNjLJdrXYdtutVq1bG7rbq/aavkCOvK
wqlM7A+8Ag1q65+9LaLJ5TBfjszKViLmnCTAvfFdy6QEb5/F10PrsvVKwvDKS7Fuownfh+/ZGWdE
y5PekBjC8YMU3lbKfZZerVR0ppkcB0nzckEA/tR0h6ssf8v/1PncQMNfOjbu18u+gbWDt83xHQm3
X2cyCQZCmLRylO9whga1y0MFOhxJ4WlmrL0rlj64TeEAqVdV8vyueUZKPQeUDxN5cdjtapaEBB+e
4N3cnRYfUfFZexXCFvmTd3Xj69jGt68p5UCAh4SuXjBbv2IFfNZ7TSubyuC6Gc3skQ5rX9Mn3mAM
2iSoi7CDdOuQri33L+lA3d77rOSs+b1OEtQciKW5uj8oDogFCSiMPM0o3luk4OM94zQPMjg9ECwb
ezrK9MeHGmPuwIHTCoGLSB1fnm/Eb75wlLnwD6eeOlvSL2n/mp6jPbFuOfgGU459m0kgKbByNS7G
E4OAwyQ8AAH6OUgKQwqvFOjG2DpwWxtZP8OP2lokhIaeGjU7X0NvcSja+tBE4ndTr8Qlt/Aqw+I1
Nd4hLJRXN9mVaq7blOad89qdQVc7bLb0apsKGii53n3W078IljgiyDIfMzjpTJmnkPTG2KmZBCcQ
SeX9Pwh3iLf9+f8016O4MGKzA9osxilgWS3hpQPVsZ3mbRLFsa8AE2fNrsD9OaJnzO5njdePQpfC
Sn7+8UqLSoM0+smRM9pbWFpTzUnb82CnbN7o4PSIJom73sm2GT+sVYV/yhMdhnuY0Mznzy+gs7NO
tgHtybqAfDehEIhzOGKVDnB1hKBZC4H8YkHzp4Ayys/oGYBSdViugUd4hBjnlo8ebJypfEtLKI9z
ziqCMt0Z78AJZtCHYlDiFdgSEK5rIPmarF6w3Jk8DTkolajB+S4qhg0HAjXfmcArhj78ZdWRz6Yz
RFVJyY+MqlQtXs4qSXJmWsvz6XDRAzYYkO7LzdlTxbnZl4/ZQe1m3fKQHWY4pWqFuC+2YZdKQPCZ
cBcPhFlw+XmQkr+0IV3oKU7D0fBC0ddO3cTiktINDhCB8aEgVzfvl641l9BMrm7U8J6cP2KeTeV8
m0YXACtblZ/tZnSkD5pRCDFrTmXHdncHo97ROVs2b4q2OHW2eJk3/xLW1oxJnLKxB/wRpNxRedgi
4/x31cuRmWDXuzQJrfJBzBO3S+fVp9vdfU6INWREMirJ1Ff5P/pqnHd02fT8ZM+7eEwIQCF8wz0I
ugEu+iC16ZroHFXC1E5Nl26UYiiza/B7DHJ02M36NW0O1zf1GGfpiNZMIuUZBME480GSdwNjCUa1
QxYUHbvxbuVXSRfFOfP8Pm5/XpMEYvMblS2knG7Hk15ccodROjh95Q/RGh5nEyYJm+b5jL+wAoSj
dITi0tw0raPdzaTnMrFrgyOBNHbB4c5izzojr68J/Auu0KXnC/ek0Bkbb/YW4s+jUSMs1DLR/xwF
4hx/qJg+B3HBPLr+ih1uUTHFMML4FJYBb9P3mgwRdmuvdjzPMwMhzR11+EmyQosPFYoNbWJePtPc
Cfsxs2l2yhlrvnflUULb4mme6X+b0qhqjkitJqtwwoXVjISysRt9ERNJxphhi+DcGsh/+o++6InH
E3rop5KgD7Tt9TUZeTO+IppVB4Te1jK8+a7Z2oY26Ox/1g5x6SYZrlJluqzbnjReO7a6szQ7NIHr
xSke5cVuMLUrAAhE2YGQs8XfW/mecprU2j5yjzWbBgRbRB+x/roFcF7Qv3rqTIrN6HnhF/I2Pr3B
iDXgEulza1waUGHfG2fTA6NQ4UNwur55pIbhkusNEITEBiHvARcqacHrVsE0dk96n7T/R05DhKKI
fpYIgKnqL0OMqUtzTZSYw7KSl4A7+AY1WtIh3en9c+ZJ8jRatQuQim+qyb5iBDBKuxDh0qKY1gc0
ghAAl030gweAUR25Xn0d9CSKL4jE6spipdQmkfv6trahj6SA6NoXCZst7GEfj1fROdJ0lRpYtYfC
MN2A6oXQ1oRWca1MsFC7rqFPU+S76I9miT39Do9LcUbrfBs/P9KQKaftz19LGuGMT4G2PxnGEfhD
4CGxtklSntOYEawVSfo14uTrjkBtPMD+uVLklBmMoOausSdaEjzsNaeag1TkIan0j3+5VbHHUlC0
aO+XRQImwX8gPgjLYnKIZAmHAkz8Tpzms7tbTbiGJ5dKVVtfV+oPnh3wXNXFmcbE9bnqIIFxwhLO
jo9rMBA5FDo52xoRW1ZQ6bNG1jSrh3JwZj/v3ROwl/5ShayvwN+R0K9iXWKvZEW200tgK1hMhUHC
YRrOy9M8BsJC78qUGywagKAm8PBYAws1bRaOLcgqvUF36JPWOrKMsx9iV9ALShS/VRMZmAFgOy4o
te4o8wXXfQHWtWIgGc/nb6qntGknas91Sy8wOPab22+aotdM/nnFEgPxJw+qMnCTsgwVz5S4TlYF
cwQDorZc+TUCX5d3tvROqMTPoVWY5htlIo0LN3plYHP1sOVNPAKpFFng2caFRQsBbSGPun/JWChM
BO81TPK3atf13wqYQssLky3iuD7fAkXMrMqAFeR/M3RgUHUytv5F5HtXTBp+/MtXPgTXo1NpWEFo
U6mcoJGEALnq6syiQQIbqOsa6XMoc9htcQshfgS5q7SuqKvtYgzyO715vDgt3mwUU3Yt3DipWAqq
10al43uC7iXNjuPeuQoZUoAyRqQdRFWhRrN3N4MZO7UzIphjQf/OvmiXNtdA8nya6npXNvfA/0pI
TYhLHj97VghSpLPUl81mJaD873pDfObtEK2SbxUtV4A5PGAKjDHQ+Mvmm4QIwdVIUXdEJL3iP5qS
722FDKaHBRneu5zd+b4L8gEmvVy8VX+MJgvQ4UOMQHZx7TJ80OHNR7F+LI1UWVI93I77kGWe2ZW0
O5ZJXHN8HTdVSWlEw6em+ALXzk8lbKXcjH5B8Fir3PflWYOUR6c68pFsdeCzvnNp/SpwyiWuSGqR
kRGDZP0pftQI0x2vNJ1fnaGsgs2GYF6mZs7D95Pw2mKAZgbcDR484W/6M8G3i5CF9a2fp/KOKKR0
jXNsFEy/WGEUXEbK8Y54V7yjJz/cx+RqQqz4eVkOWlOrE1vfqchU7CPa1IdLa5SiuCXSKW4jH4SZ
AlGZ6i6ZMTT33b74LfU8irkJJjEFqiPP1xhjKc1N/9NJXmMTK2fRFCje375wPIiexlDJrqCIkhEP
fZ2u791sgUj4Cuy7S3kLYe80SyGtXAfRcqX4WkmJMpvt2Wj+OIJ0NGIBTYCH0ZrH73H6ZMj58rHe
Rx52nyjqoLConW/8CAu/heqo+hrK+nsZWs9o8UmImeKTnLCpbBSCelD8nPV5SRd6Q6BghJ0+RkC+
bV4+krrwL9K/foR/ir0BQ+hFmREsRT8ZzZqglIBw9xFNGxWNfc157egh7ZL4bQ0Dm3OPYehnNcGc
QZNTV42VOcQxwndqAZ2Roh7N9pW3GFsRxHtjQvbfH7/+NXGOu/ZeMW1+v37LiEhHTXqoN67m6s/g
TcEsdK6JVLm8iT5h6PtO+0HenSVitNJVcP1dBo4YZm/S3HndJI+ANBmkaBBPZ4mZt59vRhppL+pS
4RE0pFCKmmRxQUsZ6ywpX+qiOkgHUgqTaOD5NmMPmU6BbcbnjN5bXZCrR2Ik1Qsyk8bKxlqWgJPJ
rZbgzhLErx8X+OjqZwa/qk9cpuNJk93OdnBZLIh1a6nmcxOg3H2/PP+c+FddLf1axXwDIo/u3XOW
mBFP2GZkLRHKqS4MabTrcumqQUmyaw/YQvWTf3m7CLEpeiWacaKsnW5/SPc756YyT6h6eQ1jNriF
dPDeYtWTmnexeFmTiN3NilUMDEOuGyz6HkKElFVwCSBmRgEUht+WxPmbsaVn5le07W7mRtFDWTYN
YCi+WmrnpcT9oEa7ETAfQTJ+VmtJ0aGV80u0z2mAq9hkO9bRsB42Z8d2m01zApd3niBZ6PHhuCjx
ZltglDY4LPJQ+WwVZeP700mYkmMthQElEsA1Xs0lyohkf4v0XRbel+9nCwqmTdJO39CXrnJjVRFr
0/7mW0vw/xgveOY0I3CczKnRhqSj898sKF+PUpsWzytM8LpnoKwO113C/i4xH/xc8sEnSw2Dsj7m
yq/kq1DI4g32rTUbIMauf95jiyvRAxHO34B311pcNFnupX0arteQ8TNHSBq8FSMz+20QSxxtjiM/
nQgF7sVWcs+Zj5fje5xONGaVwwx23LsmfpcxNnVd1NGg2vNDQFiRt0iQSnSg38QKpm0Z83kqCtab
lVKsxcIz0ViySl6EaiEqBN2FNPPlWBgp+55vNvGDbKrEOVeerxn7t8gkN5nJA6zYzstkAJpqephS
TzX9Vv5PCYlHxiizUPK7YbtxFrIBk5n3aVy3L3wWeRFVkIFVG/oI3cDLQqvGxsgHfhZn14S/1v6r
Y/khJdaKv/iUT7CEDxQDybyAWQfebWFBC951FXQcUpxHdFPqml/owG/uSd4lpcE/pspqgsVkzS4b
MzxPrgpGQyQPWePY6tTauryJaT1CdFlF0iA8IKlCUlAcAaE8ZNiBisXE29mvFqO5iwDoAUcSXwUU
vAo2k3Gl9XRvnwcULR0vp1RxcrWYJShi13MuOOaJRMqMxCRHsInp9L0ehyoL4Fn2/uBpGcEIpyhf
D2U2Q1WXJwpm8wCJ7/UTPcBHvSnYGoMusTrfQs33trH0ox2lWOyQj/pQ5eU9j1RA8rJiWLva2PY4
UvEUuUkxf3sPk4QxnYZLO44oLg3681bD/AxXL7qYQIhG+jAX2dALDxJzeOFlfDlIiwRHnrHz9U79
zQOMt1rPSae829pVbk3YeZPVj3UcTbomUtv2qD94feer8STat1lWs5bZ7Ll9iyOaB5/9XWLH7t+9
3vp/lmyIShgeNuxIrAQ3POIQb8EzW/4r7iWXRs9dxiXtfbLYHOMb2MH6TnV+P0+TuGCSMrwxC9ee
DLQQhK2NyAmY4WgRFTQ94H1gbJSS5lRsbYvTAvTnF7nnnBjWc47QEHk6yCuOZQ3mxpMGDkCdk4OI
AIk6T86dDBd/hO8sH9yDrgPGHxdnmFuR5kNSy9lZNWLqxRNf1ZSjQpP2oTFCKDp+PavfUD1RPZX3
hBEJpsKKo0JG53EsDwzxo5uh/59mvh99R8hfSAtotlAoVedQUt5XhMVdH8pJj84pI0je20UC+DJ9
ZSEmqOGZhi6vQwVwSiRwoMR1QPF/PNy+0QvKCPeFJMu76THFzAIF0H2olA8EAcl+rtu44Ncvvqg0
92Mo+FrR1vDdGZ8xeQg7OqKqFakEmpSbaHWxUMgHw72K0v6E13wRROFl0YsAqSumGLQy2g+HV//k
DjJmH1Z9X5XEftE7DJtC+LaUXGOa6N/s7xirguj0h0+DS5ak3kWEn/sVrzZXLcwrd8ZI2jM5NvVi
+Y8S291D7fNa+W9Qib2cN3CYT+/bTdsU10o6t40oU9umcdNFjqW7OVOwJ2C/TLMyjo/t7lzpQR1K
X01okBVommoQalQjGZ07AP1mDvfisxMUQmmcu8fleMWruwmuRDcMZv5SY0mdCqyurOALfLnMRf8/
dITNmXF7nGtLoorC+ps6pMo2IauIJMwTe0EgM22clORlFnz3eJTSW298oK8OYWK5HlsPVFp8TFJd
R40ZZ/brIJSAiYGGSi0+ivzP+DoNF1JnbbceTclaF64YcHPBnFnAStbJ9ppwHjegw6xBOxe6GFVq
AUDuSowF0ODfe1qnihVa4hAaUFwwWq/aLMwFOxL0oOXdTgVU03vJTCadPFgX3GhCppvypqhPlE0v
hR2pmaxPtqL8IFSoocgK7yHgtcCVGR3OwJGstf/TuiwA6ujSXc1dYNgNeNPuQ3lYhKZ89JAOouPQ
TcCcjaQRfenz4lKGhXVzM2vXY8uQiGitu8jhjzi4FIBF9EA+cE1cXIgKj4DSfj+EQXyMPWqT5m5z
rRfPtJcmiw7tbmAxKStpzkHAQRJuONz/resbmKr5QYUVsINdCOa1Cv5Um8k+nw3MMT2XXhZ0kjT6
QH00RD5Vzw1HQZ3kZz5I1PrMqddQP7LLNihInU8tTOD7iidxF/DGqlic7YWOX+sGN9X1LEYecumQ
nH3s1dhprSMHJb16runyv40aFT1voeHVXIVoPo8Mz9muw+NWDPvX/x0ukCsmEd6Vk2oCIDSGUo9g
fuTM1icNnwkTfzbG+MntpRnGX+bxIDEFNnJxty1bWHbxMrDCvtHqI/4Djmk0LwnikHpoZcX2pFrD
UqEKx+x18jWVl4YArvJkZbH5cE2AVMiPr1NZRiUeeG/nuD+C/EdUls6XVogsqpQj3Inj0mHQw99N
Grr5LKBPVWW0htXTk6wLp9EfD0P+oHbVIyiVkDImNvpBeAxDRTyh8jlA1nzE8cZ/i2FIfxSi9YmC
1jgfs54idfiOXaXAkCuMJWSdU7gGN54s+NsNRHaQg7MJINOT4/Fgkl7z5ydym8N05zdnfvM4GZNE
w41UjsiQp8q0O1bC85NJJ7aLSh9f6yZkU++eY3r+tQSlItJB+4Ssew91UkU3tvPkKH3YJv58DKSk
DIyOKNhQwj44vdmM15LkyWaOTnD/skTRP8UGiVjNzQMvv7KpGxmRVMK1pKd26wPdS+THcJ9D+73V
Q83+C+lluuRgEhTfJZYRjFEh0Fsnl3tGRFa6vwhegHk7GRj66/moVDB5Wrd7qmvvVh0tVcMe03yk
GQ1SHkga83ILsneSorzDeLNa+AcTNx/N7wfbowYHwVyelt+Ij/cWAjk8SVMIn/xjhpNSBmnIcAXw
jJD5ZlkO1e+pnceMlvURetMJQwpWR8e6ecyXvaYaGP9zi5EZ6RgzodSc6uRi1vsozSda18jzE9DL
/eCQHlDVhh/SjCDHT4TPZ8xzrEVDpI4e/hqrV39vGPpJHFEMfb//YdzJZFDXLooMZsrbjvYMBd+f
WBhqRdqe6jooCvFLhr8kk2JJc/lR+qnHWjhzO0kDm/QZgiVnzL7CEKuI64gsO8k2jcmsmaEMEHjH
m4EQJW7k69y2oaQNqzTx1dZqjJYvXt/eQFjWZ2ngjPlQjuwWsQxT3Q+Ts9i17ZQRjjs/mKrqKrRr
Zcfn3Kwp0Zuu1b6P/uY64wpTGDhS5UBeyQMiMBDaqncH9J8oCuO8OsJPUvKGFxREYpUCJlQOOON2
E+yv6J0Ff09ERZuzBHjqbVTETjucOCYVYz9ZvkLtODSjE7jIAA6csqldI8pvHloNHZx5k8FZbQU2
2aQu80/es6kEGSJSOHvm7oMBhS0zKPdgDO30XDEaCTyscHpmVnoLuyB4tIHZID9th4LZOFzxQK/w
XdIsndVHhPMhMcXA0SnSIqygwMxhEtCtMRmDbYtRtUQZGrvNOXvjpDdayPBMbJUdeEm3gexjOlsX
+KDeFsO8ncE9tAJjB0VbxSd6Yf/QnJOCuMyVNrvJTCZ1ehIYopZ30/fOh0+NUM02CfbJP7AH2KuH
ABFcSIZQINsT7bbfBJWZT9D5g3cpSppmezquC/OYOQo0idyPGwLsOmIoz/cdDrotVamlr214m6aM
06+P1kn/TzaUIRoJXkLxJDlhBuo90sr0cKgwVARyYJvZG/awF4Ec5vthCZlrYzpqjWXH4ZDs/1Ea
VP02pv5ONnR+Yverl1boNg/kCFqjke69ddQN41q2VqicQ1QYPVoLqDWteL7bK+1Hfr80j4ebCTB+
Lkf5kLRYnFTOkA9bJRuVskleNjXSslkFI5s4O28q/qsK9gLMq9LIxIZYs7LIDxtlT6QPy3NMx2ws
2QQ/l7pM3XoOJNZ/c7q+xAFCWwhg6hMujlzYGNUrEtFhfkE/r+/AgsQersmI+GwWfxVrtz/ovQqi
UMIKGFplD58rU8sBpZhesquFc7vo3eO8GRhYYAf+JTavRUFb9PtF2yF0jjikrmO9p0VQbQs0yfjz
wxMQqPsnMYHyYAuS17qDrdMcomLDwiucTklytqqbFpYaUTaR2tSXSv7InG8oAa/r8IzZnrVCfEFf
0Le48P6iOj+qFZIDzgSjvCVaCZsocZTrjj/qMoqlkWOA2Wx78AhBZHRrhp93CyDCilVtNGjs8LqF
PBxfiiVxddIdSnFhAURAaYs+9mZYCSMosPx9J4ns2QhsYNJEeUPAOB+5uQDMcCCeRCdv+hnwILyZ
mFrpIoNq7B9C4dXQit0POxjAY6m5fQBXz3QCBOS+CM371I5JOfoviu91ciw3o5ek/fI/p7zlCxQj
idbYie/7e2sE1dPOExHNLP//oXa6XnLsQ4G7J/UWjKBXDPT9Ys7hEmCIy1WdbSephwUC50WudU5Y
gdBbqrjUbLRqZJch35ZHUwkOpoZfK/8FS7xlh8k+4D+zFT35S+VcaV6R93rwKN0ZwQOp0+GLNbgc
jxs5fGwpiXtVI5BzitlqonFS6FDpVwq81YO2uMJXdhX+++c+Mxt1kOrcbOJTyBfxNiwPMjHg3zMg
AOxGXUsWoZcROkPTThOSfcrvLQZhctS0oBv6+IKArB5VAJXGrpwzATAAD1T8cm4d4ofHhDEtR5j6
Bf9/MOYYwKFKafpzGbfBE3uR93MxJRT1+YjshJ0diBBjZFkATqI/2IfeX3ElfwW0K63eT5mNWEgE
f2KNL9ySCBzkp6VaBS/30uGmmD3obNDxpclPwydfD++DOFcs7IbaergPKegq70BO4dQqg4vG/yZh
3T9RizhxNBhRej8GePBLxNRDym93QJX0zWz/ICEqpziijiAD+gupejKXJX6RJdTLr44eN5+HL5jV
WuTXteeXomUyaQJEle2Vmm+WXiDpjQlomf1heZ4Jb0Yp2fhHQF9Foda/Ozs8jdFPeyHXfcZvFkl5
zBXAAQLkVAdG/wTjE3bXdfaxSbqDJC+CSq4mRk3IYEAF9A50LqVHGP6FhDKLZKonUpaY7rsEzC2e
2fCet/5s90oiLzXfYFgPKTp+JWUtuKRX/tlvNZznpTWfZTICspAMMhDzJMcd26N/QMz+zsongbqI
BWPXcp5wVnVLbkQLkydNbxVVACq/OAudD5mV6SN8duBxzSmrowq+ZnTttQ8hkuNIVD0beMNwh8SM
zOEC+T2IH4wLFhEmm5Fo5YjDvxQQWGrrcRxWViPFRyXNbQejthOKixh32hAFQxRdn/dpQSzwDIPy
yRKjqk8uPzE2Kc5OtUXJTyC0CtoVLa6DbUTGb3U/d5EhFA/nphx/W2af7sJP9eXO21nEz/M+dyDQ
eMsqvomN8aSWPFG+U/41m/I0hgYxyXF90Q4N9uXRTyat1dJM+YyFehnm4MLASZVkn3F5UTqYGTHk
tXd9oHQQCVPS4fZhOwV0H8gYLHF+nc5P2WrvjCMDmU+fY2Doj1PKd1j8RyQo02vGNIi22o+r6H4+
1SwPAw4R5FHcC/b/kFg90PxU+NH7lS2ZNTmwZRew7d8V05reJwICqrsq2CtJnqNPF9gt0WVTaKNf
kbNYp4LcPgIeeIKU5acvYrDEO7tfLCfC5mKCZjxCyvGmLCxOUc76+3+6389YDYqerW3G0A3ZvS3z
xNSIMUU5sUenzFyqojCTsalUjOF3JzCBuZPMMT8oy/+hHtcD9lNbGhHMQQAqG3TZrFGu7vax3XBr
y4LKwXC6eV0I0K3uR7Oz5P/7K+YyuC9kR2SwERXjgXILDzDvxgaxSALy7V914yIouESrbUA0cmo+
56tWqILpBKVs5V2l8hZtT07aNoW5GxEZMN4MsKqi/hvQgXYDQGejA8VAfr++gqpxDQYWlm18BsIg
t9dnYEJQWwvTtCbWJ33kRz+8pC7bROcVRQ8DjwIx5D8A64XNHI5Z/5Qp9Rfwj2OghndBR8EwSHH7
fTozieNKKgVVt5AmjnoFjsNs8Y8LmP3VohkvKRtWu+YFgtjpW/gZsCIMFNLdGO4gaaQldNWDjCCl
Kek8vF43tgEkNGYyZPO0FvZeeNPokgJNp+Gc9mlpATXolnd5E46It6oUCCvcCAN3hva9QfZBIh7b
QyOp2TUdHBX/048pPKgdfJdwpT1NF5aNoFmQJWPdjJniWeAJay7oYnRfjxceIUuq8zblyJ4m9094
AbjnFVPrZWPTe7klHw4jnhjD5JKTo7wqwnSZFG3dWq4G5G820oAx6cbeQFBPDYBEiOfd0LkLTWdN
88m/l6QtTv1u18Ro+jrB5sqlf4Mqm5oDbuqUAZtEfohfenE/NDTt3LYAZ/rzubWjqQDPKjYYu1yR
pjXVcJaovL0JJsMOvUA5Hy9vjaE+fRKyk6ApzUEpASZ6FN35N5GEsG1+9NfGqfP/c+H1KHsrPhP2
iUSW/7NCIMdq3pzDHiQAXbPHSf7lR1LGa1BLdQ8Njpc0W83NCwwlhdA1a5vETuaox+Va5Yin3LF5
0IiyrlA2S/JSJkRX86B1ddEK/pAvXT1soMvPkajGQb3rpagXXtIjb0pxUd4HEJiBrZfH52GqK/Wo
DjoHXpkYisAc2w0ZY06fhe6l/UzCnq4EOErQSX7Tz0Sp/L9AURBqmdtUw68ViYfwhni6U5jB3O5a
LOVoOZMjdLGz1ycILqfRDSi9yyl+Y2uARTDPM4NWm/av2zVuEj5KuI/jJ+QOx67AV0bXkO30kNrx
cycfdrT1HVh+qOen5EjEPdJm0YhXPGTQdGOn51oxmt4DduIOizLg+46pgxgBQnv5iRXI1B+5TR0i
0YD6nUJLgOnwNP6qRaCm6zy750U4JsQ79Xebbjtg3TB4kvyaCiVR7Vpzsg2NQtHdRTnuVYhmGWAt
PMvkEZYCYoqTGLbmRhrHDwx8JuxdFKObufakyNE6AeVhqX5uyU8YT9g5RaBxlwZ1kkLmBE/Hgr7F
sgq6SIhYFuMW+bNvZxYQWDXCAODUOPv57xgmNoW+JjoDDeQu7URP/1qadSjBMAJqrzGtQXr0Hn/f
9zErDb61z6OhbS7TTNI5sGlOIkgmJr1kucHxeyMZz44/qnS/tCUbxOjDeIckq7TgN/TP0Sy/sZDR
hiLIsoyR3mZmxKlCf5oFHeGR1ogs0RW1yHOp1xVHvbKSSMUyUzyvzHQ4dgSDpkzdFihBmSJKwlKS
SfgsUDI4Wby4dWBJVuj+ubz7e4Kg4XmhQjlHVz2XgVE85lqKHVjPYfixnbasUODxJZOs+hzZ8GzR
OaEfCdYJjly3vb3fX+IQsaax0goKZBhZfm/DvLBXq5nSj+2q8VLMMvCGvZnDffgagqZkrIhmpz9v
nUNkFcco5N15TS87wGg/kMj7gKXynhafLsbgwT6X9mh7udLP+lwjIogQ4gALZu970raZHaujgVUm
esago0wROUTAF+nfu9AH4JsM1O0WBc9wPlbzgP9kMVboXcCncj08Zg9BhyJlzGcfc5CxIZDtJvrb
N7x+LO/BOySp8WsS/pu5ymmgywOyQOkJcHfe0Z5Zsu/9AWjYpCQtNRWDN9ngkj+t3VPFeP8Y/ZTY
4aVg93h1lPz3b8KD/OIpvthclkilHzKSMaIxKrCbefvUqNpJvqFSiz70svqnYsvckMsyKmj0uV5o
+Z93B/Z8ucAV3zZ3aQjXZNyI39nb/vLVUa6/8TMH/jwV6xNPlLFrXgicbdp1j9y8h7g4j2TPuMIc
JCMX++C524xbodWRVzN8PfIAYOR0Sq5JVrd7rk1g0/5IsO7ts9khUs8Sq92VSEJPKCNHLD3hxZO6
Szuril+vSMVOFlNCpYxiVxA8c1CB1yoPTm167+vrMb3hrVMGPz88zA5XsEIvWX4UDJrYzd6wsGVO
9J6CSNoG575Cn4A5+cfhS62r7p4dEj69MzD2kQyrd76PEEJD/8rAQVFxpDV4R1X/uR25al7zwMpT
MhF52pQiTnZjXjH/Np9D1uP8m5Yjlmww3m4p4ZTtcttY3zzFsY8vOQEEiKyhA4dWGbXOiznUVx5w
QlTCwcFG/RJIIf1+oJVmftLWoYAu14zV9WCSoqjuG0h17r1MOkR13CHrxsQNJbfux8VLKIrd0ybU
iQ8dtpQiM6xVWbOTi+wsnM/IGTgtHbslap9FStP5eL3JvliWwcc2+9aCslqIxarj4IO0k7FsIAKv
brknnnWxuT2TH++znsoaWXlRyqyKZi3t8GipW70cU3vTiCAlFru3x+WGAgmK0jOurKCtDGx5vpx7
Dsc0hDKrIBj47cElAcwr1Rmb6/OKOLeJsWKI0AwGKwk11ELjfChSmwLpWyT7jm5xLyksoTRFYDcA
E2OOPsj76wY1t2vsoKM2gCjcqzVLCSN+NNUU26ZNkv5Mw+uBuXYswlB5mmwlHJjQVPR99zVLbwvd
5tWAzgbRUik61ioB5JJrYF7v9LyiwVXqzVp7+pnQVBGdgGI+zd4Ym18Qh9/dKi5Xc3Udo+k0cN8B
Gax/r/VNNWpDnEY+slvu7strBQAT1erfizUxaeA7jSepNKNbU+GVy7DUf+gm9A+fn0TjCwCxZgl4
WxXJkrHVKv2wdH0GGNF0KKihJuKnXGzx9HbfuxHpeSya35OPZCwB64hRi5JWd+X61ldjjTnY/zRi
8ZO+FtM6JSfzkXKhKozyEMsjvCpg1m5t/nKQJHSeQhrLHmMhHEdqeFU1swcOrlIcs5ygt35qU1KP
OKylF8/JjYJ4kFZg3fs9MNGhyHSbu5pkHYizriFtSOPyRTNrjGSZy29VUlzxovwM9vAurHYcCe4J
2eVctWXxCqd6uDE3m6NAyLWCDz3sS1zYY9BWqUxttBpU/00w68DHPwfsQ6Q/KK37t8meRWj6763H
bkofsMV7vozER+zr5Crz9tAWnEEQuJpKjsJNvn5vDmNsZGkocszZJ5gdudTW+H195ht6W56noZq9
OiAxFU0zEzv7Qmn7ZhcrKpUu4eiRE8vD0jnqsDxnZoG4mhkMptYtuaVQXapfRn4sD4tIAvFomrvf
v69iQhwYQc2MGiq5BuFVILbqf6tp/cIlsfhmp/n10B/AzpjNNXpCTJA/49I9i07nf7dtOle3LuW2
0fgx/MmzaQUkm3Ua3GjogtBHk/FIYEDiiZjaJor3bv5HmbJQbK7HF1xpgbd3SQ0QNuTfGhh0OTnk
HdHZEX0lm2hxu7bpwbugjSKp7Va/wsukNkeDGqT+/GqHUDVZ9aWam1F/I8WIB3dlneBR/LuA9RMd
nnjPoOZqn4XbAl9TJxS2FrabFD/GxU7u73Qu8o6vkszTzDJJhCrGMAT+v4l44TL5ap0+i6caZfKS
ttW0O2cOcSQCi7vDrWPjLC7WUW4BWF5abnsH6fRNJ51zxKHjeiO1ZxjX1PxGJuUZDQgdZjsXiw0B
kpOfXO//fswFSRVMhyO5/RE63igE6+HDd67J8EIQHN49E1mVCqJgo8wrmBoSgFMYQ1Yj5SHLU3CM
ohiZctKRTrFoYhXqbYW5O8qlVHUzZtZFo6wFSiEJlyYjhtf8gQZO/Dmc8GiFX/vg4K30CY3EsbHK
5gBkBreav2cZ73At2zlx4XP63Ro0eLT0ZZagXbJzy4yN+mzaPTyliTpMZrbiC5/m4/d61Vz1BaPX
p/wjpWOAoAu1s/aVzbBz7SJyfI/eOpGD0mAjrevLjLlTGNWHXD3i6CeDsxl3IDvLVruBvsl1c49/
HfYo61OHyXt3v1F0VbeuHc/sd8bI1PSvJ1W2Gx+eIUdqTDqq9g0o0rqoKEhooCgikLTeY6kT/rx0
QJQ1jO8xnnF/Tcp/RMtkH4imBJCkGorelelEfyaybGvi+1yuu2Bj/N32y6T2kmwS3zpYuPs6R5wa
2TIY++FjjRDYGPoHH0z2BhJgZDNi+7tR8BYlUAA0Vpm1K43KoGXy9kCNbH1PrshubcDqlNAqffuN
REBxEO3Ju3JnGC+jWWxkbfgNIylLgskbeCOe89SOWXFE6PvXVzNbkWG9qPbUDPcYx7CMOspYs478
7VvhXfBdGzOrCllzXZNADubJaubdMtkLFjFDLIREPp3xzRJNDzac+kUYXmQPTR/Sss0tGF4L+50X
nTV5BQZDho8G6ADJoKscXwJa30XQG8hiHufbMN8AL4LdNDXGD5N61YxYV62/xOM3EZuvbneEPov8
iD+qaQADltjF1MP3TzY+eSlQxW1pCKsSc5C6RIL9kaClA+iMB/AsROCa81QGMdOASraj+tTUIe8J
4G1rgjgGoRtKpRu8QeFUS8+eDr+NsqIt336BP0d04zVuAvrdO50fjFdRqlxNUdZpFnddEwsQFOw6
QJ0Vd4RiBMrRLRhuMNjuMyx1ebLeGLbZcnA+aWhRlfbla+xG1BI/me+c5XnlOB8/chpMczDSYBSd
o0GxqnSD+LvdD1+4m4zJKlc7wTL4hyCMIfE/TEqZo1GpG+VMcaX2nHfSWN8CbactuU7fZGEHPXk8
ceunpOCj5+L4B5sHFjIrC2YSMKMrEyourh3b2r4wZwWRKVy9CpV9ZDnWvFhGBfKq03LuhKlkTM6u
+NzHg4b5OsqemWTtjCYFntZvu4P6kpuNf2DZ8rlWsh8G9vqI2xJb62e3tGHhaSETOtUmL0C78Y5j
HSI3guGRAK3dNIO5xKWA+zcBDg+EQ81XirjyPQgVuPKvd+AjxAoV0OHxj72OC9TOCjueRwwmnkIE
V8aCBdbn1ChaUIOMXVjPW605XYm1XFaOvWlcAYsVKGwpSepsWacHFHLxQOsQXNWfko4MW30qdKZv
0KDJjHw1iav2mYC04VOCBJ19HE1Vl5uWq1ul4dOOpc030HggPt5PTOaU86P3XbhI8lFmn5efUANL
PvvOGcm/wdzE57mVb1U51hkJzy+VCjwliXwb+GdQYAxk5bH7WpL3IndP6qiV7//Ps9WjDnBRq/Ep
YtZgIe2jIIbZm7SC9qNHmNQsIuXtIL7ZcLEHXXjIoMAEeTXdLolQDWY3Of/qTr9ip/94vRml5IzV
R9+HfaZcZoKAD7tQylj8+QZOJtaQQiqyQBdb9MLvC4S1TbShZLx5NN81Ij4/K1IehFHTus/QsvWv
OA2HfrGwFVouKfqWrL+qupJpMyp+b4PsAN4QLvMdD2yTCr+OPQMtPwM3SBVsqBpA8FF6S2RU6PQj
L+yzB9fMyHq+8buoOBNwcYAH6aPy+QYA6S6iAHLS//W66MVzsi5eQzHmyMfjv7WRT6OonzvZ56ME
qvCG1XltwRW3iomMKT3DoqOjch4ZvAIvJyHNAwvYhNvWzH2R8q4o0EBd0DH2TVBaLll9YCfA5q7E
Be2QmfogAqJXn57KD/NgmMPtBy4ylkTRcIeShIZyR5Bhhiu2AwMST0m5eTOtxai8zbE0q7DCAjLW
Rzbo4nA3NUi78RHpPGjBR8Gc+J3j9KFuZ6vdwGde15o/8om+PuEnhBCLHMbKLt+zEnmljpUD2a+C
8JZgHjORiiNBEqQnQOGTqP0LfEZb/kv+8PCQATQzp51ke1NcIXB31lT5iZ0Ijw8uZey1vHyZsAid
j3jnyuT+acUIIqjCRfZddo7fqZkWxEARzPfvYrUKBHEwyEJlpDoW8jVrK07OQGwRMM83BgOXX7hF
xVK6kBwHOWG5YlK1OIqiMO2HIK6gbA1P2GfDpB5HG5nNXL3tVoo++SQhf567npoWLDICns6KdD5k
Lm4XlUL4XhuhJCDXuBdz2kmb6APd3aOxlWWKAyDrj0GBJLLj7DzPkAwSgzewNnvIUBN4g7VgEKVa
oR4gkyU1eRoib58wHsH3WK7JPmVPymBWIVStj0Ph/BrTO0e/UAdCi6ZpkoHYCUSlbINjWGjcSweR
HmtiPw1bPIIH8zlQvRR7sKNuEQDoxWoaHNEbrkUFNmA3O30kQdfx5Rqk6x9Vgh0kRYFdGz8/PJiu
HZaY9guhIjh1cDs7o8gUfwhEQjN0QZwbsXEi1Jx1N9NGK8aIzhwZRBi7gNNehjzd5raiNaqJd5jA
2Q3Pho6vRgZflwBamjUIc3TNsOPoNWAiRRH44hdpjrNt+ovzQ9c+PUwUbp40P6tfg/X8GdXIxTG0
LvKrmBT6Py5b3rFE148gwR+fiFpFEGAv8s7Lgl1zi3MzHrRXKcrNS0lOPwLgiq8F2GTN2jFgjwPb
lRkjVZf2jbS4DsAgyUes5jvROcvqHakDpyNm26OpnMPvQC4cViqoVwNSAamTbUiriZDMUuzyeoF6
rh5x82W2qDySKRz4F9GT7ZR0X3LwRw8aeUGHdAODarv7JLK2am0YFbEo3qLeJLQfJIONNnxtPj09
PprhyMzASfTlayd9lbwoe3DnaB3ws2802qaNBZZyLw/Tl2zrol5qtA28tKA+gZ3r3w1IV+kl8xiD
CaVWwU0CbjTlc9ddjvnSTskrEJE1Ozo0lnZDX3+8X/qSthXF9aM4ghgh3uL6t5+2Rj7lpaDT1PVV
0FDRQd6zPYL9wDNTTYWKi7kLjOKGMxUKXDf7InB4AWdB9yvUHKcQFYwuKmYj5L2vKI70124YntDU
NxR/9kNLlYRv37TjagziXSSJv8EC6WT04UhYJlVhXYvsWBp58wg39/jEqpaTRFlwXjfwsv4ZCMYm
+2tNJRw9E8yw9WsXRfMmDakYYykSjdiZ2fKZVDLwuJ8Btu5mNQcPiYXxzYJUPsva/kDxkHPvVezj
59ZDov+8DX9Q4iPjl94KNhxouXoFWfuCst+cvwTkkgNA+8X/wN5oTMPd9q4b2OXxLolxShwSjckq
jeeag1RCzCX1GUlP9ZmRXkaoOMXXQJP37RDoKILN9+l3kJSRr/Wp4lBqpvjeG1d4RRPI/R0AD84L
3qXyTjjPofu9mAvnNqExMD1S2IhezMWwfZznPze3BGDWJM6daS6R8vX0bGD3BD7pIfjPbsSWmBRC
uUA3Vi8J3ufO2jX75Gq01ZJBHhC2TlG8NwaEioNQKAbNVbE4wz85TT8qfZoaQjVP9vWeZfaDOPgV
Sc06bDFkC/eAqOohUyTJglv9/nPRaswJxPVZuGseDGgo4AKf5+ku1KVluzZx9PYaIOV8f+LEBbIK
/R4bRKCqgphsDGyXnO7eyhVD/kt3YGxEKBoJM6Yubn9ca+yPHzXwnirBT3qcV19Ue1jeX5hopw/T
4jHrk1Zy+J2IsiD4k1nJXj673d/QuQAALyIehGUd2FQFtQyiuB5oRgjUvB19DA4geE+wlyApvHk2
HwwGKr9UsTw+D/AMA6SuGvl/yk49OHiiK7rej27HzP5B5zow/sPzX4qa4DfxWPK+PxjKC1jZClMp
gB+VTCSJKc2Dr7JboDqsx3eBt5Gug6G3nek1L7Z7cVB3gVFrLeGh6qjhQSQXURbfjW5tArItAaDy
RxNYo311B8/mYdmbBW/dYAqjnWc8PH/rHZDDumwAOTrKsy4g/1eUrZHu96Hfvpr9gxvgGs1iwWFh
8ugc6nhV+penoFV5kU/37bKMG+hY4y6a66oQn8kDFBglzaFnHqqDsMojqGZKZUQGJvXPlQ1QQx9l
HG25LfxQcSUJgNZFoMb4k2tLFDWPJi8qSh8YizRutvNQU75X2BII8EwrZx7wKjr0J3QzjgtYV1U2
wcTjhZjek97Dqn+20N1PIbD6lh2zUmR+229yf5CODWyZF8UFy7Vj6wJX4BzF5eK1GI0npEtPo8dv
QsIAdh0qccNtK/LdsTLCKlKAtVeSlWe0B+wrZBdKEbUgaUJfp+PuBub1Nkf4UwUNrFNmRaLsuMAM
QT4P76sQZDfz0wAl3Mzm48Cs12bjvjJgaNBZKuSvk2049E6vrKRbgTiWe6xkp48eGdTpqh8TDOeQ
O7rOXhNVv9mdQp5s9AtoPI8wGfZaXKGRSsaw3m3S88szHfXMd0Itx18wYAf9f/TMB71ybHWFcrZP
Ymz5216VrUzSu3Ba2cFPQjspJ68pqjjV+PIFBWPr+EXIuBAzJaiZXp+f6ZDMITL3XLMKN6uPjZmh
mVxiwz77n2so7YjMPefntmq0KmEoJvlBK9mBTrqUMeO8hLg3oSV3Usckyu2aW2cEdTfRytmqmFUx
cLHvXSHk4HvPLMlllgAni+4JGIsKKzmhr/7gZAyOG8vGMDlxN9//7GZx0kBuBHXfxAsPTm6s5HFl
PGWBOjDcC6/eikqcHj5V+WdNvcJzqNhko9WnyYOsLUBUEciIAfJrV842OwsICgsHtsRNZKgpZsS9
ygSHYYTHGF0e6af/Jr3chLZatfVM6Fn2CSG8lHEUABC30JPBxqMIX7yYjbZRVHed2j/hWG0AN6DW
Y+Oe6gMjTYLfgK/TjkajdgmObGSSrEfDaPeXtZmypekiAd5c/obBQAOJyTiLrzl5JTU2EjaXLUES
nAENfizaTkIIxjw4uM5W3FfiaPGwQbkTUnH3MWnqjFrSvXVQ7ODizbrWSxTDQQgQUn1PBj8Td9g+
ymv56dqCQYh7hmdbwvo7a5kppvjfbXEDKh3jkHbTqjL0gT3433aPWIHPJxLtHt/KtADjAhomsiRY
3iHQl7KWLJkV5PcbgTfrS+/H+YD2GwHmE9uf79PcFXWog7VMFAVOQGlOEz98EJOSoZV71FOMAIRB
DgPYpfW1EfViekkA6hDHDTxKc8Ga+X11qQ5i7DcAjA6YKTbQ1oyZe9x1UZW2xJIRgiI3jwmeZ/K3
XQLuH0u5MJv0GET945ogwGDKIzuhDyqcareMKK1cKZqzP6khl3kQ+4xQdyTuoATV4c4ZH7CS3151
6Rz0mEc3qwIXX3x085UPq4RvrUMawobOJYMUoLgyYicV+zfrwtM09KH1lp+Ri33UdODaN8RyloAP
+kU1zyXVOR588xmt3vCoqN7BRFavGoB7y2PvNxgLzIjl0Ep9ld1OyxWdeag2fTioKyRruzkRiPgU
0bx2qvUJgPkn9OQPW5rXsTkA9x4VpSKNdJHgg1IkkVIxh7uw/pjDst8ZhUGo5Y0tKpQZ7/mSWcL9
a4yluiMLddGPOBDTUFR4C+uzviVmjbhiTwkFR1gNpywqG80Grvl/0gkHqpDk+4wm026ZREx9smBH
KqCE38Edrr76TTvfnZLbROlpLxdvdw0xrFg+iUlL/7E4PhAWuIcOj2cLi0gYlCU9ad5gDGJntQ77
91+caYxmU+L2tv4f0F0lRux08Y93+PKlfr+0KBkucTedLaQCE9cqoLmMWP0xkN7oWcfu7BKPvbvX
3uEXdJLrOIJh5xHeOTS+aura2W6i1ky7rOkb3Zqd6iuqb/CJfIQ3qA2qO4HKqoyDqVnplSnGNxmd
GxkDROlCpm3SSrsPjrNtfQzn3UAPCG13Veuethkub0fIYtTDfClj2zV0ZzRhpyk7ZmX0ecdb5va+
r5d2JIDhUEWpNNwTZtSTpYumbopatNbrgCxlq2BA5O8+GaOWCXsX4Bljh+e5utaCmSt6URvq3BKG
MFKQ2L/OrkFJiK1GT75mIr9SHVkINgAMN192EM5dOzpKDSFtcEZ3lAlamScjCXu/jOoLSGlT1ooZ
yTGaU5k209UjGIRowaoS7kawOcVu35t10wmkqK70zokqLIGXATE/CnMID3/MEOwGOEXRoLAtH9xd
42KTlzkKLBU0yRRSL/tnw2OMSqVsN+PeN7U265sWO5GL6PARI5n3CNJXiasiJWO5XAlmJ6uGN0U5
prk8RH7eGItESBWQEoV/5K+zxT9QRQfNUEoVHizMy3ZP1d11jJYVYgTUQlkEe+HD9lktCqb+FVRq
UXWaP0RL5kFi4ATdZG83WzIz0SObMCHW1p+l4J3I0/rO4lfoyOxB+rLT3+QsmPbKWNwekEXduNbq
Y8GgmxEAHDBBp+/91EqNpYg5eDtPyU73asoHwduPRJMfvzwmwubXH0gshkjQB1QeMkf8NK49VODF
iI2zpILKb82kRvhR/UcRGWYV6F8PCb2cv8NqaEfUEFA8JQO/xA19mbnziYPLERg5RwTAvxqBfYXt
DvImpEl2dVy1auQpKR0r25zgaXAgQcPVbGhd/TkOKjbjS5aJS5ZsuEiMnSsEkCe86z82hGdbxZE9
hR7iwydyS3pw/KZ3kj6jaXC8JfVcClQkNbm71E52a2vjjUw4TXxgAnOjXjpHeOlqbHrRdSClyV4E
bwR/IhY5qivtBuGNXdfnbcmjgtMlbe6HZqmbHwneqG805nlrUQoEVGzSa+Bz/7gBSc8EfRmxQWHr
xJSt9a2rPzd384KZyNxIAnkWqSCTH8+JPR2id8WbpnigPHlpPI/yQrv5RWgD3cKbfPki0p54bDTV
EUyeGeLR6seWmnG7/saewg1wM07HhH1IU/rKWkVbG9eAYb+yGOz1nUuZMgmLJo/StIkVmQWCuTiC
6tI057/B7iPeW/QGmw4k3Q7XXfIoERq/muZhud1A9X+eLJJa4jp7MzSJOTydFJQ0/fzak4gtFSe0
2Wr718ujD0TSuKIPW26tS/MHQu8ts29HYCoK8QAi9n2LY+6xjxrLRG3GkXvI43JZDyrfw1U/7n7A
LiGZZPRrMOhJb+aiJ5iIfJ/ohAY28RhsiX/GzlZLof1Leht9VYuYg9G/YVRaoSeKp+HloM9sab2l
gnKs0AptFoAnuEhV0o8VeNQXx2Zoz9O+ZTT+MASaDoIh89XfGc8oc0ecQxQIT7EZFJ7GfOe8vxSO
jF3QrylK5+P+J1SIj/qZE35xB9lRSWkQA3VhkL7A9UJJrth8b4FScTdz2Uxv9+eEuWF0bzf2GMxr
d1f5gwn7VXkd1yqGs4LHwo8qfphRczQ2mupNA5+/5/BuPt4TNpjllxzAi8ruPhwttj9dmp9PTCRx
LX23p/r5gSYLZAnF0RXmBV3OLKy8ifH6CET4Hh1YI2I5SCemn41zCNkM50o1mFxLNbHxJLjr0jWj
Rgm/R88RA4W6I7NpOLfd1D9evr6P2P6wz5iNo8sVyQ91aFe6+HVEVI+tNzuZKxQ+eQXhpx/p/z+I
3SZfnxX91wnGJ4YYSod3XhROif3EhZ05Nu5b7zE+wlm2mC7W5WHhnWMZxLq6rLTKZWxMaz07Xq+P
vRsnxDiLksWVyz0n7XOJmzyhZoqU+zeApGYISORD1D2MC8HY5cY+NSAwLUBikTTK/zfmXF+sOluI
ob8aAd5CJnHD8ROb0oVj8C6fUxTes1/aASl+ADj+6zuMNb4rmtZ/75ghvMVov53Xdor4bHstX07H
2F0fhUT8VZesWsHsRr6MjlFRMYjHv4BCvNBacBfGPvc91y3L+hvz97yC7xvzQ/W8MD/abnOMa3YZ
zD/JcLI/gZB1PGs3Z714ieb3D/iNiBuvspp6rh2YGaBbgoibrcSJzWrgfDj3ZvYmiacKRJxRA/Hu
AgdpY6pPvjKpNeD4FQoH9/noKU+D7WLJ3j2hcL1TuPLqCRgShxfKRHANEN1aYtAZScSzbQAC8MAp
O2IZ29PV7yheVBdMa9nTr5MIQbzso73f+oZuJMbqUIzTFnD7v9e+dNR0VDTvF4G06ncPHFm1PM6U
3GbkicYEKnmO11IjDkFqhgt7tMOeGRyT/mkDPVBYrkREGDhzuEXGGVMITNM0jYttMTSASBEqpmtQ
mDO+rseMdU5+FoaBtjCRvf219c9SMLMomhO4i5xVyCO/TkmcQzptzErdexIsao6OvZjlAOWgOYns
EuRB6XYiNWdQe6pFK4nFuy/LcayV50kIjuAx1fhChbbgjfXjGORn0QPl9HB5duD76PpkZaPHYhjv
wesiRqrqZ1ixK27l4qtvgAL4q+LiyvjEDGW4BoH+xZRXmUlGm/R+ftjWvKQd/Cqlze6MY8hzAdMz
hJwKf3Hik+7kvO8Sf/rrzSVTe979OIl6iQY7p2TzaW7DnK2LujocDk/FkK8q9SXWddsJQDKhm3vr
dzLciNKL15Ki53mNDzpTwoX8LTQSnK4ara8v/5+GUnQ+uw/22Zqbi+QY1D2vQ4ZilhuRKKlskrff
bXEn0Zwym+PVTGuL7E+c45sOhrRQYWV1kCsrxAmwGlyL/S8NudrgGDFv5lG5B0cstwun/8M1AUgO
ANJvxvxtBVNiNeaTzK+gMal2aUI5RmbCr7lDPvsHaPenaGUgmiwowyhAdzJrtBnTueW6l3EkBGdl
yPY1uvRCBgjxjlOl2s93vE6siVYszEXWDywtzh76UiJhnBnRAPjF/jCVFJPOcqYUulQ48QQakD5u
SGD+ebqR6uWNcM1wNB6mbc28Y+aPwh2rzgfJ04DpBvGjGazC6ritVg8ltDYB/jbd96Tb0YlDtmFZ
033jNzgz2ByrBaHYfLGD6TejvAw4ZU159p/Egx7wIH9mVAmPMaPrKh03TcDOKaVnvyGNN5TSonj4
DXei5YFSOAbyo/vCpYYPtPnLIxAIVyUdTTSaEqaI6Lz/EJ9eOV5u+80sQiF9X/p5G+S9gnMjztfZ
PyxEU6qKuYoFWl8qRJdkEl/909AOnzCerUEXjZ4MVx0RzSj9R1z5ZzQocdk5HBDs+bSadGHy2nWd
qcydRszaKDfCUkbfnxLtdFRZuDz9revowN5MV1M6PzhHTg1BEwujAm5J/X+kiX4vFg7AAsAdmBsc
ofsmDMD3reoJ5tBI+L9vdlnftiVjkgQUEb+u/QpWOsVZ6CpJPn6477pZ1DJNH2EFMZBIFZlevBFD
uX86MlsCgVok2s+VHtsJZNs6F/vF2Ec0AE7l9fsJ1o9Avhy6ORan1CrktTz50Iguui7BRO4hE6Fr
BlKjuF+a2NXPRpxdLeV7d0Fm8AHGK8b1r5xmRUDHZaJm29u2IZFLsbWhx419Y1Ntd779Nb0jv11G
nDa1HuJ4GK3FqgJbzh/1upJK8Pzm7E9z+8OoN3/3Gq0vm0eiIEoebNCGg1czNVAm23Kt6y0MykVF
sasNLjkhivXsqxLBdrlClLbVOviZbrK9I9Im1k4ZxaQPnf/u0rb7Gk565dNJyX043wr/C++NBrSd
1O6iURdiKtfGACYiIUp4tcedQjyMy0Q3RCRhMjc4R0Nr0mOTcuLZ2De0KQ6ciMrUnkONbUEZy//r
zlyd1eHtKRthjYHwGNltEG8UgtWs3K5G44JYd9W0jgTuRrD7detVMMZiXOpctZ2YaA8YMQSHYmtI
aC1M8zny595fk/oS/AILrM8UTGTAwI4y321WbBvqz8TDxmllExfXDqKv3y7CheocR+mxO09L+6hW
XHf1byOhNYr1aat6rnUvMTeHXEQtBqk9dmgT/8m5eO5aI3+rn3CBa/xOLmZs5Cn0BY68GXKP3Ftp
qyXGbMHhHkW7XbETb4b19OnnwzJpGGQoMUiLzHkMXwv1aWlpj9BNmA+XKxNx9HyyCHTP8xOkR6IL
p6tyGk1M8hmr42W1RWSWirIVBmz0PAe09f91VF6h1vvVupOzOh0YAytXAVRrs9Uln3djwBjZAbMD
PgHDvN/PXMd/5oywcZ1gckd/oV9U6+U0Ct49AtPAzS5DYUp4AAVQRwK54O+d3b9eeRtB03mKVRRP
ejvtj6yhw+ovyz6kOWAdhQPODkRZ/MDqjuy6eS2ya8sVfh5s3QmP9hYvoUhzpVkua9zjKLKGoo31
dP6keUKnW+DoeO6XGMldNDwX0zg1aPhCRJazpZSiJxeBh2zKi3SMl3jH9LLFUBsg419cIUii+LrN
bFFIA+4D+6Rw2SlsCbM9ftsBi9QgpNo1uP/9fuVpHfL3G4D9xNdBwog7YzSd2q8q0QCw/x/a2TtW
m1vwkzuAKeF30mW0nBc2Y82caU813UqKG8Y7w8S+CiTpSzymTl2d7u9uADzm96kE3o599noDHyJp
QgtVg828YrQqCqIh/rZZpDElPOZwQuJKjSuctsZAZGfRTGnfCh6OMDiU1CSZ0IhLjlGaItEW1GU+
174HWzcBQeAEvNN0p8RTAHF2c5VegWDXQdc5xYcm+4IelmY+5yZGorXmwcL9CtWfUIvHkHss8Avj
bBCElOiBEv4U93EqS+7LHB2WWYh75BYKCTyDnnVwp606i8qrOnePxW/v+gTT7K+pyj0unGacL61x
4BqLYDZNDRGPIBKz776K1mu7yVRMPhx7pysWwLceMYdrPsml1jLC1w6KlHrna/iDKMNFVHatFbfY
OE7M9jT+Torug8CMFLy0Xuj7bSZDGihQBsqyUth22dxny9IgNUyfqfwKf6Fi7o3vOgGO2dRb1lkT
1WE1yGMBmO/nPE4oXMdFZ9BBlhrbzCW/HWkjlMhh99QP1dDTWZLIcAOZUEO6ps0jLyfUN4GEcUdY
cwX7JqSymsoOI2K7sYAOv9EHb7dpLaCRIKPa9W3KAp1N6YNnrpDHmM7C6hfqN10moPU18e+clfgf
GPH/XI3ZsC8rxIXFynZBRRiTSUaG5PhVZwD9eUVvqzei8oeiYAZjEA0XjOokqu2g0Cw3ryfcHGC8
AN5pNjPuxfXVe6oFX5XDM561wwPXBP2Ldg34PLEgiS7HAizqabkcwKbffvzPmKKJXyAQEScPKqec
gdZCK3lzhDDRheJM1WDlFrvu7he2DRcug08hJ59S1lkq7qtepAKrllND0ndq2DXGFeIxoH4inkiw
JPQzk9AJVMXBAlBcvRMQrc9R1CJA4pmKelc5jfRCvf2DIiG6Sac8qicPL/sNtX+SWsay3YjAaV5r
6Q7Wf7BOsi+aMyzVlvYpIj+CSsgfzPEqreYJ0rmEluVPWPR6w5SI6iUtJ5Gh/O9E4xMZtDIORKNC
HrssiWCPd9618ZMFhJfzIT7B0Hy46zAaBg9yViKgllcleVFV/cJLEiwIdXP/vFpKsCIJbQNzSSnc
3YH4SyKkv3VKNy7K7a9oAMYY2XFRA9Ly73/HSB4Ohpme3uX6l/Xq5I1yobyExbn+E9talKjIvR07
Rt6CiinvyHgkPGrXZS6WDb0MZqLmcegwuv0i/jOUVPXeHFjVqf4QP8sk0H4jP6uukwhkgUzdYVcf
SiX4Di+tSIOvp6ohSHjAoKo4tbR9ZwJjKfRc2W2BfpFlutB1lLpT+Ws1KCJxVlVOzS1+BWP9JRQA
yQySsnhp68+JIIdoFnmdkRyBn5PygTede6MrYsqhvahaOFuaklrOgOGL2GCjgXPQSWnrS0nIKDhk
wW6HKU5HX2Pt/d2ZsUZfmkRpwfGRkLCa3S/mTIKzYY8MHNNo+tM98xTBBiAgh/M4FW8X6twyXBFz
UAeRmx521Idn8NGGQzcHNlNSmmtAAPNjjGyrfrxxe+GObOT1BryOqoEQW0OQzLy47AcZ6lGPEwuT
FIJUuSyyOkBk6DxL9IavINusMFmmc5bQEOd5TAzf9EzyoJwBsLb+WpFXiQrKuT4RnihaqzLw2H7p
79kLU4ZT694rnWuOAbSR+hc8ifpsz4yT3bveEFnRSaXHHDo8np/QKm//9NPNSEPGOCPbjo7v3EN7
sl1Gf4Ms9qVCyYJjWZdrSvP4P/XeWi3/qEGvxqJ4X6rz0yVSikV79EvWxMbB/z1RGs7XJWg8vRpg
0X1ECYPLqvDY709EeTtBYycpqip73+5kkSyDMY1ghy/5ACMfkFVzjTFg/+1qWEnnuf+NeHZJ6HCN
7JWb2Om4mr6jG/qtu4hvfCIateDDyBub2xSirBA2tGvAfEfoCr95+dbwd2+7wKj7N5/jDAAsyu7u
lvXoxjFVMcJmFhofpLE9/mav+3hctXiIM98HvqnNThmjRdaoiXoz7Mn9U+Ktx/S8duEWcnHN5qMF
UGN9cctX+D3BRPp0BgnoduCZi5SxbZfF3h+KMJQksDk+YBjtvd40AEqRoyP5JejVDzLwaBRMBW5u
GzbKiFxKkZFogcMH9q/T8CKoW1aabagn0gN9bMd6d98qh1FjX92VHuoahRR1N37H60/Vc9xQ/Qhu
n4/qOJZephkn+Dz3DbcMPPt9fkqKFiK4t+p2qAmWUvh1GgFUUqRXgLpnQ5w7YNkUZzqa6k59qDIp
ItllPBwCJw7QM4XFrm7VeAJOzVggSLCASDPYwJiMlPz/fteu9LmSy2JCnPWp1leMitdPWSBzU6Qn
RApOJVmC2vwmD+SrOnsuV/qVpnRrqP4IxAsmQx1Sw9jrgvPtIlK5Jg3MpemwPAC1TEPQ/M5p0wsf
LA7GwPtNq38TEYMDU90D0cLOlQOczbuAbMxx6wDX4N2fkvu8I5HZUhKF0GUjbPkLh+5M8BPXR5w9
8T0uWfNNFXQCyM8thHp0EbdULoG6j+l/nRCj04gzOMGlPSiEcbuhnfV8+VyRCpVXgP7fhtEZPYix
71kjxCXR+610dP97g3/ONYY/KuKATdZitSJJMogcYVJMvzdDp/qQRziFqcGI4BNbhB0iky7hb7mx
XvAxOnt3Hca5yzGEqBTS/as3n0vzUa3TRfoG7Fw9adzku2uVACgX5rgYfrRYWquwnoLo3V+el1IS
BBOICbfkOjDw1nTIy6ljjW2s+VB6XgwTJTfWdUPs/c93mszCLUfwltrddTNIm+lpUHuRAVpyzfxG
m6xvxzYLpXUI1tvoORrwYpLIifPu53VMODy2SYM32bCZyK0CCP95aoHwO4CtqSAg27rBzK6Q1T5Z
1KZBKdwqwEX0Rn8ol1h0D4T2RyddFnUVWNIlRU+Laabi+NbkkOeJvE4NPaWnsE7e9ZOFRXKxYEnn
XMt1WUNHRK2IvViDQElukO1aeg2oBNW+Lvx4fecZ/e/bMyHuNZiulxE1ti0pic3rfM2BFKRLeerO
JhdbGTMSJBBov6BFEynY6sftRfUhrh2Atkw0aPsDfB8shSe6MJktLS0RgIqFPse2trTusjlWys/n
av3xwHuSdBvygELQ2R0mqs6yIpV7041fewAcTLmhGVZwRYTfPHw5iLR35jlphDcGGT3dOltUDy1q
qyiPNi3TTYTJiI4JXumn1K8wUgSPqs6zXrfI+QFx9iXb3eBrUXU14M1N0GNXOsu6QC6HiZeMMaDe
vy87c+iaXDC+/I2pmLLkCx6bMeqK7tV9DirtN+KjtTBclLXXTCTLAcIzCu/dI72CMbgaGBUBDOtk
jSQzARg/zRQTVV4gULYQiV9DMwm/Vx4MTxNetJsaKCfDibDG90tuw3+9jbmTnQW9uVgxI8wzy/Lm
q8Hiv666YjkaGEUaw4aEI6MakEOuWg3yVqSEqPjTslIDG7JeOVpReQDFh+/Bj4Aqa/WQfOTS2atk
IHbEM0/1j6/bBic1dP7rRS6isXJv5AJvBJiiXoKDB35ZTlokHOi11pywmDJ/CwJcF1E0aTmzIyUs
59aXne0adeA5cGmogErVK/NLrcPjdP7vbejMaYq4BsvFb56SQAvSYnxC6l0+WPo5KzfYx+ZxwO5g
ayNA6K0GERCVzYUCihAmsxx/+O+pAQ9qdwQtdlDSTqXOC8W67A0xIf4g6O4ILOGh3JPSMU9d2F5S
CASgpRH4RcrBT8I91XEWa7xCf3MnMLD5zOrUUIK5HsnqRVp2lfZwi/TH+fNBG7pDYs213KhSOMHw
Ye05k+Fc2XxEemc1gKavN3+14BJ/smbLT3697b6mj0IS7ezuODPGiJ/ZVgGh8uha0/SSWGAIx3Qy
hWn1KJ8luQEkW9VK/wo6JFBjF71pIezdLgWxqAk/VlSdPcl7beEYVk/w7zvbPKCYpTigKC9ulL62
27V09wScfxH+DmDSsFXb/cOUPQUIxsp3fYyJwWg15ugH3ckknYakBfsqonnBtkO3PbpWG7I33hQ4
8bvF7wE+vwJLHWPrRsrNRFd/E0UX47aIH+eF6x8nmJW8OOU8cItDrBaHuklH3/Mm6SG1E0g8SqcG
AGZb/PaESkm7TxhRtKd/wpSWR71VEg9hpSrMmpEw8CrfHDPtAvnq7NlJokGjww6pHAAVraETX8s/
pkc1CtXnVmlbMxfCkA23Ja+Fpd0Sir+zw2p8VEdX0iONT901zfyzEP5CMFlxM9MYW2Pj5RAXbkMC
IHpCzKRZa+/6/hWiRZPfIpehbMAyYyPbo5ydVXZh7A73Vgn7zvIWi83O7BFxj+DVqFexgcUwlQ8O
Mbfktg513c4e41F5CXcQKfCK6eofKeQw2vdxI5hV+aj6rDDslohM2UQ7LuJ19pGMr4+CNC+stl+Y
AFS9ZZDzIKGYAfLH9lGVZT77q0wUDJEr+qcGaQ2LgWhyyWuQt5eq2CAPiW8vNu3PCULqPy3TnPe9
lxsKAUJFm3T4zsuYgHoOssbOr0fe7XO3ErFd4LZMqwGCp/T6ODOr8r0BMJH3/7mzJUUKUC+QM+R1
/fY+6JBZkBZ4U+NhHgqqo61N7NBQ2bREMjDyrzI6V4+gpHlMQltEBSFSgWsmKzJnLOC27bCQStJh
xkURUSGNQXGsnFYwP8GQ5twvVzeg7Llk0lYLEC+lsjgjsiLhLB2erYbWNr3v1GWcY3n1VnXL43zY
08LV+CLqhzjmHUEqd66A2pq9YgcJqr2RqukfctiBsuGY3NfDfBopQ1EevPs0YBnb4eilkqD13UJq
Bekw7SRI+kgdlaV2KGwmMCV+LcCONSE1Su3Omv3KK3CDttlw/LXPnsrZ33Web4VlfrQCmIF+PxJK
VkpkLUhLRwOvaP63sDZWq9Ia8lgnyUbgEF5M3dJwuZF2nQTYbsvwOiteT3rV3V4c4wh7pFFSVMcx
wQXjgSVGb96QCDP8XL1iFbkqgacek7oZKzoEqty4vry0MuVNBqNtaCagwj1EbCZJwDLI9FU2XoWv
H/0l6ddaGdF6a5ts0vOq7dUTmahW7AHm7birq6nz0XW6PRPV0F5OK2mdIXJ6QX9/2idw1OvgQ+rB
R43Qgd0lc9JnBpuk14A+3cKqpnqt9MkAPcXVBjAkc1YAIb1YdGr/weJWqwWnSigmDICqXNU80ORu
VFgh9XaoB6vJgkkxRXDeDx8G6XBvOvHoKvpkOjqn6/1Wb+ddkiHbWQDfp+5sT+KcOtBnj7MPKWKH
5Blz2bRRiNmLqbElxKdiUFOarf4NNLaoyXCysoHfTaH2cs9xF2gmywQwIvlobQjkaZhw786HWy/r
5RGqrVA5K0fbIbbiVrRBAnlqfQS7LmUB2eHUEVgpwKGo70YDXdgR1C7Kxc4jcWWpXrmXg8ezBtyR
0Q16ejmjzjdbURn6bAPM464BEd8PXF8EqzTzDw17l2gBBQwVD8sCsszCy7E/38d6ny1+r01gK4Il
ZRJdMr0Eaqconl7hix1bQbDv7qaztcrrk9xfGqtzk2bkMhFVpJb8VHO/Zik7tgRTlJEfLf3jwiu6
WO3UkyhqlgnOIrkf4UzU26o5kqYEjdHNqNr/1GOziIiaBAe6HfiubqGSmtr6kPpoxvwdAFByA2bH
iIR9r0Vd9G2rcZ3Vz1+9AatTsh+oEPzJSLPitjMZKoo2bJ0CCxlvjp92CUOuJmF+ZzojBD2HPwL1
MXSASo/pRYn8m3r6G3Nw3zbIenDZV40zAFAu6e4hc88o5tiLK8u+9N4PbMSJuQO/xsF4VMoNzd+g
AcgBO5oJPdDXq6qssx+AM2KTW0dv6ULZ2Dy5nEidglKgkehNBpZM3VhNjKZ0HSxyr5m4+mn96dCj
RIjTBvZPd6HVLwx6qSdsJn7187sbLcIU4IuHEz4mtFHfy9Qw65J4gkVs386ZQz0/s3OIkK4DL/jJ
6q7nAaGp8H2IWxQAWhMBkmq4gKmYTs0ivZDjGJqQqCQ6xnjQcbfbhKkvn+NMF72AnTgqzi4ST1o1
ai6E29GYA4MSpGXf78KBSFzScEyZsTJV5o7vwwZz0eOHrlaBAq4MsUj9ZTwD4H4Fs97LIoQMr5cA
gWng7K5TBXAKJjl2hpfb8dnUnXYqzk4mUk+jwqHr4Q4gm/52j/wznTVqvzhQ670FPY1zWxRqrKkC
vmDbaWwichnK8jrYUj+mk2MoKXTTma9Z2nmqbB+Bos83gySUanhCKp3rYyVuhabRNvKU2yqeP/Ju
HnBJZUk973izwrZrfBqcFp2JEq/wUESXohgULAxdPgQmIFYGLeyXggxdYQA5Cuy31iys9fsn3chQ
ssbEyS/MwklrOQ9UUMHWUZuCmXRc7mCmjFuUY57DpT9lyKCDVtdwYSc9cCePomBLVua+y2q5/+mU
ppWiXlgrdDkagTG2FgyeiGlcTlLXtTXS5jwPbXbQqfsfjKU1wSJ96SC5Msp3csr8hT53+N1pNyXY
N2DqzfOkgNSYOua6zibRCjve8hWNIUF6RYCuvFQ/4OpmV72u9K4Wkdp5vNHh17HsMDf2oe/AyR+g
tx9Du6qiSmqLMchpySLAWe7d9dcjlHQRio5pp4Clxxhp8/BeFC8yDAGicygwWr+I8U2b5o6f5/Ed
8rOKx+Hfu0kQdItCg3sPZJFZAbwuHyuLZU9FARWuhoprfE4Oc/drCW5AdBfVocYfOH6ktpXNd1cf
xKxQhYR4XZrZr0ONDBtIobkUUaOu1ONKglZgVzd4fwtOBbbOzuNgmanyNVoCYD722ESagAaMzODA
Btr8YNDzbJkWWpagxtK3ma+yf35D6BC3wnL1z6EkSXcrp0vreYl2U1Zhkbz5hzmIYajE2Wj9mwVg
TqLkHwDmrW8ZwcFlYZPgOHxBTBwtT41TjOv9rlUi9bXgRH1K9OishyN+5GyeDplHHTebARDD+Bfb
RQnS7lK9SdFZSzqn1x8+UFSQoSJRpqIcU/L/7OjzWTmARi6/CUNeO3tP0iINikx9Jjx51LmgW3Hg
fvZmTG9jQ3JFHexaQokwSNflcZmjyVc6qXbpioS+uGZZFIPpVNHSI/Ip6+7GrfHoezIAVywCEzE9
ORG/nu9DCKxFtnM92CQHHozAEnKBmMArLR1IPgKu1KeXDXpfdmahI0LL0VMnmJfxt58+CaC0JgYH
l+su9s+OfXxl8kyCoOSn9z8eTdd9oiWb6EqbQ+YI5hCIxlhd2/WdtABHEAa0S5MdEzXN61c4hi3i
2sFHwQXHHoPfpM1e7VZGULHADCRnyPQGL4UZp0yCOfUzi5qgARdLbTgCoVJvcqEfS0B8ca2rrlXd
SicqiBkYUeFvafgj3v5nIxaRIAUTIEazVJbvZfLfD58tpt3V7O+6s/eW6mXkOEUPGVrC2uN2QxkQ
YzO/8C0i0aSMNe5y5G0As3R/48QK3x/GA3MM43YgS/j/wWOAFkCALU1NZADMc9t01x3eCzZvX2qj
LBD+GZCgfB8LgEJe63PBjrmBOyc3cMSqlwML4WL2TR/9olQ4kY9+/CbouozFRZFwui0a1Y0bYw4/
n2FbfkIN4xCNcPmp5dRGsMxFFADe2evIgtZlDWCiqnREvmAlC6rU+xFV7t5Qt5GtcRM5LZyqMxPt
kPp7MNSYu+ayiKYSr1pwzZQYgZQ9B8DHoN9OwecIXW4l4utM86u71xqz8FzJF6IEb1NZi5gvFq8k
3ccGhitrrQytX6zN18eyitLohKIsQRyF+auMQ99LlYiX/9Odgq7ObfHNndM+I5kpCLHpQFI1L8zO
bXo87zylMCt1OCmkWTone6ifpYxJX1Qn6QVQ2km7XzC2dW/jub07sLTa+71amZPtqvNW15aixgxv
dPo4vk2bZw6ZBehQNqFrYr5Xtda5ASorojonJsmfT/1En0IAIZLaOCvi9LuZ67XVecEUQ7wVHc4r
ErFB2zSuBzRZpuAr9s+364IeAvDr0/nQEQVRHYhjk/AUbqaw34KkDYgxYjcfGbmQNL3FvQU21fGe
wSXbfREv34QbOemSohbRJiNQImkyHdkOxGV+mq0ctyxOw9yR33S9UTTKg7A5O8hsitsbZNIpCj1u
UNSfGuq7yLzdG/m/1tHRDAEXGcKboag1sAL9jYDKGQiaip1D+xVwi0NaKTSqlRyfFGEE039onOaV
wPNHmSIUDTvLsAcqCwaVozhEWGnUaBrIUhLJl59wrpcXeTk6jnpxsjvT2K5xL1v+QQ8td2bmsbgM
q76dIvCGvw3PTw6zV2+iTo2ebSCY3z7DQYdmCV0VIIy4gucq1zUEgbpB9ghIqdprmue1nJIErn4k
7OkCFRyLzeh1dyFSuRwUCKHZhbPddJzAOEBhRflz1cJUIYV88kW9idjPiBl8NXgYKKpDGMIh42DE
zIZh6+JHAMtqJT2OuiezJuClDs7hhmCaDWEa4iWzcBAWxgaJ5UeK/jVxyXomKSclr5wbTmLAnIPx
LtIf5fwcKrn2QhjxqCfhs1Lqg0h0Ifiz2yQI53f3hBOvYX+h23LE+/wyYVdwuz7/YHYCs8Dc7uPa
A+fjpyJCVeZFyNGXhjXs/aElD3mTSLamMyMED6Sr7GgngANmiKf/WreVa0YV0lDlCrIATcEmExKr
Y7zOnjnZqHq8MsRlN/8okRA9X8cBMCr/2VA5jrtq5eRPvyE3ShlHI+pDlxBLL3/k2iRPSDfH+kL3
EIKQ+1mJimm3FC3TrHey6U1NPo4dckzHTUmBBEKjxrb6sdquXXWTEbk82HCP7kb+kuqaNrpCd+9I
KuQ18hZ99DOsucxlcKEOPt4hS9ReL4JiewPG/a4AIGNDkxygP4wE/wwbrxlmvIzwKBA1oaJf/60b
w63wtJbgz5oO8nxjSIowoaSm8plGUDgPSEurOcsZnslK1lGrr3N2+ReOUbe5lP/8jqqyD7Uyh90t
IAA5VJoN1JuMG2aUiqL4ASHPd+v6ClYzIbHNGAnkjSiY3IuHsOIoUxqRkX+nBlPWC4C9YiBI4VLc
V2atDlJtMWGu/jPNdo+slzcL6Sf6E7wOQznx0o/DdwqmkSYO9WMlAja954A1xYOsyXd6M7D9Xezu
Cs1lkjM7AfNMokt8vRI31i8OVTUGXgXHIS86DQR++t/avOJQOw5IKMZUmPDKVl4kIKtFm9hLkens
GKYIzCbzAZU64gkDxCrfwVAFRzcz9uYraT+ENUzQ9y8o+gZ7Yr7ovb3ns4Trd0Ybx0nYY43JKQOp
EpInfpxfxm05ANbVIasu1U7FxSMuKAPY5Mb0PXKJpHO6mNHnNd3E0QQ8sFncYV/6G5vQILD2kF+q
k2TGIEPjPJukBnWdCTSe3TClgguu4fmhde59sPvEyFnpBODSZxT/mxnqpA85WKniv9qP6eOSfnDU
dfB5/zr1/eAzfZtE5t397tn35HKmxMcxnfGbiGfD5mRfuEvtnSpRD9pdfOLRgqaFs1BbAczZjGBQ
Z3o1ds0gUFShKMwvc6YXr+g/83NcH4Z9X+sF6tHkraOv4NejzPy2TJBTuGM54oLvW0OrlWsk19mI
u2zxCBRfxXOjIw8evHRo9hNx54pcdQetGEq7eLbYcHe1SpmVSd9YlQuYeEG6AZuzNEoGAEWKoroM
14AH7tPDRM4N1y/i9m4DASFyJQoPUQqyueMi9ebxGoSnooTEX2wa8VRDqSOvFaaUMqlVlaRvZRxO
bR0JAuxKP7cQggPsmmcyQXGCsR40v4eyoKV3Ud9RBqkFAoygfRaguWr0/sLdjq0uz/0uuMiRjVW+
prc6YOKyVOpBItZGjDEtfBdWeYJxpxibzEZXLkCRwg/sAfwajyh2hV0Ve+wcYK8QDPbwQVUdLLY7
oBN4yhVI2rwj5wxAsi5Tf1lffO90Tpzytw2rcNWxaO6EaoWoRo3OY2SKLzqgeLFP9VstgJB4GpZT
d6eg2qRoL0onhdhKeihnml+5PWj+bao9d/tXDuaVUT8n911EcOuLFloSLX8mJkjCp0WqdnnUYb+v
Urt7rSEDiYzAxbEBmvGwkpclRALXmwykK0coVtXNJ5E/TywQtW8kRcolYD3LpYvuI2ehx15SQKf9
XNMAMHHaQZwZzq/OO86fkbQOdFTDptmEutOgPLT5/QSXj8QB6xvCBQVIWyZ3Yeb/PXX+AdZZaLhm
9GXtg/kOQfJ+rqKxsy0FCtZn8r5uSx8rwsJ9m2pNk75HHtlwAVwE8uvGh79QeeaeEukykybQh2cn
8B8TRZulCsr7+U/XyjdJiCmvM63u8iGCdU4L1UjhE2ByTCTUl/Jwtr+dy3IrCApyEqd6lxn8TKL0
nvuzYvgLF3yBBK1ZF9T33ebHcnT0xRnnMxDyuMvAnGj2YlVmUGsnXXLKYbjU4RlexX38iHzI3433
rwHUxuNE9/HpfHx8sWx8U6TzzjEQ7aIb61rjExAxMk/vWo0GWYtTNTmcd5D518Xd7n/vzfnL29IM
rBPi8q3DElmI1o7RTVSsyLGwDxE2z7pisEcax+u/Z+pij6dZ8oBneLB9KTZEtsVlYCc2rqoPveA+
KIPFl25c7NqhUaVd8brjcDJCFFRLfQoqdn8WRxPvmDPwvdwXk7NdYRx4U/jDHrUJ9+0jaNcFn+Os
CB2WyRoX+liyyZInpxY9x2bddYH2RraKqIeWvc3NOPfaayv++xi/ynjuXc3uWieFkRThyFx21KZM
o9vFWKPm3cIsWRLhMRxEMYmYqHpwj0CORnjTs/V5yKTpumRiQ4aYzwyrDnxxoli38prUuPMG5HqT
mg0P99rYxFIicoIVU9bH6WyAuOOvLbG415yxVX+1VqxIznY7Jy9oPKZnXRxLZKyd1HeGx87J+Xeo
1jF0O+nhoCYNTTBaRNNoSfrZzQWVh1D1GXRHIkw1Ea1KIsz50FO8eBiBumtKbp6naeUL6R+GIPsz
2w0nsZHtmqai8pahk2WfLloRfB/oECjZ0AN+XUp4NfHdfp9KRKC307Z2y1IY58KnM5pZnGiedqj8
h/GSdgOJIo0l6JzzgJbimGU++XPCHCkH3zUiwfnn9p2VfVCp5ru4cac7CWLWHpaTMJjZHQitSdzN
u/dQYYdvHJaCn2fzVFOyhntM5e5zTH2+GCcsSMYBieHSraXdMkDhfNEkDKjz6sbz/EFQ/6lUbwA3
/xX0OQeOw4Hg9kcbY8H/QioMpLazLzO4N/AQzdSkUasfhtYQeAcQL00T9coZcs6QdqB+fG5a6Sd1
8UbdLzUKZkKP5JHULbLdCm24MmnvjhnNk7EGRq6ZyV/+vJ8Dafg52cdhbVwMlwR24CMT69v6trra
tMVDtEkeGN9XTWPaBKq4b/g570gNwoNdTLJ7hsjaupNpAG/3aZfJ6uZEvAZmW0VTzQbptUg7pgeX
OD2f6qiEflpiRYGpXsUoLCAUuNRab0vaXLSI7tKoV79J6Jy6aKHFRKqOrmoPjm7cKvVunkuXIMj8
8me1nuNdwGnC0LPeP6uTlf6J6YiFd+CpydS19YAHjWjDfiZWmYeLWl/vVYm3ezolo/V4RO2SJ1Q/
iq79a3ySgzgina2iRSrBJ69na+4ejMLls1Bd3BoUfmf5o6kmEeqyysJ0YobmoOjdlQmPSeAKuUU4
8q8jcdJCS/KkluetWO6ldB2R/h3Y5xpM6ONNkI+IK6Ks58yDnJSCHqBn36ryWJ3A+qu9OOO3XmH3
rDEjxHf+0homqhlJZgWhCFZBm49R8xi+H1fvoS/oi5c84agsYncx75WH1J6ZOuwNhwM+Y1XiQp4K
dZEW/3aTs/npeRSbHfrc7ZgPqQuMHRvUYqBoLWzdKDh7s+BoYSFboVhL13lIn7qaVN1z9+6aavcw
elnb1387ECBoW6ankqNIQ5DFxb6/4s5JPAiZhEL9Lo1OkP30uW4naLxz3SFq3NFiYvwXy8DgNplV
EFgOO8+/eBECkh2vXarlipXc636Z3Jf6Bg/oHSFlcliCCRj2ndXdzDA6REtxFVga2Y8s7z/F/jYR
AFPRkN7x76J5qB9l6gqKVui1iIPaPbzjBayWmUPgBwOEzHXbqF7cQkJsvL2BQmRVu1aVQSm0ekUK
mkNoxYtXH+YjA29zT2GX2btqZZB3lwDIcUXoERU+W3ZlI2AEYhTSw2cSV4EIE1OG0QWY7RWKZm98
h2FLZOCp/M4KFJYDhsWaHvvddiBbOTQ1BR/V6epjmYaOw915VHEdtR0/WSvBqtnlM3oVlj0B4wkY
lHsfaGrD7IgJdxaOgYu/NAdBs8gfBXXtc/zOSIRkeXCiy3G43er/q3QNSrbDAxh5eFeHhYSjx1uW
oi0yMY9/B8CYyTsszcqiVTBERIhuMWMrqSEJ1LyGKb9cUSzEHZGRSzbW6wUpG/6QjP4YF54sE+vQ
jUeDjpO/iGCDFDby2d4Lm7i60bcICz+LcaErCa7Ua4caA6OsEMn357qNPZ7ebtBwwHTZ5PLNaAAY
btBRb+Xv4gTiYm79GNWdow6qKvbwFhsSoAvxl8Zkwk7cg9/lDytkp3CN7aVM7WiieqekAfAhfroa
iXS2XaFRDaw1mfbdtCABFqeQ5TpltCPm9NkyBNh5WmrHUohzcrYNNi+ZZSJLARb3r1N4v/KfjtId
4gtpZd7Zakt4tLg03v+ZwZZdl03J5d7EJw3p3O7hYCiB43wFm7zGeOhgDu5pzNKdga9MbXh3SzsM
l0Rm0BuDHPcL1zcvzkvO0HROKvI3gkdKQEPqTlH04BKEmrKsFLr+7GB8c2GKxT1Dq01B4xzqQv0b
qNXikEap0+jMwIUBKjnMhGOam2vWs7ZLhC5NK/7ja/VjwXN3Su5jt2SOPEa67RZ4igQ2d6psMT0T
RoDdz2tgGTScLjZ/MEYFKfppRD457WwFolwHldZFFjzxvZxvgHSX8BDxVbMTsXWaum1ZRkumcZiq
mj2mu64OnOSY/qKg1TsqpvFiZoIM93ObdRNywgDlkEZ7bZOoJe6lXYVtN+ryyiJ8fT1mf/MvhuAr
DPi6OmuGxQmpXl8p+8gPJbwUo0CmX+1uOIH19K83FmWGX0xFp2hs41osX9dNLaoKiKOqfWxPonaL
/ppyrip7qIA6jo56xEoODbtTcf5vevqs63i4R6wmavxbIGeJqQlmuGKl0IeHFlo4vY+nzsLdx94N
j+BEf79biCKNY15j7f0bv2G2rpYLIedc6P6zUXFJorcgeLXQAFmi0fyXyUM0aPVu4oseM6vK5N9P
318qrOg+VU/G96JUoD1XSXPE5lvcbOSa+51UWcW2dM1J/VP3Ho4roSnH512IsnzG6+4d5OqWJRAg
9eqMb4oCpHjW5HZB8vOT4PBTNAxpzVy70ot0t01HuEuWEeUIFyRt1ZR2BIW1sS6UX6YM3nxHKP2Z
qIjKTM21hd7XHVxu+B+BK2yBP2SxzPaCWlkYfhSzduABCiRIz25oK/NAfx/vxTVPriS2CuPi4z6w
NMi/KJ77e2EVBqlTM1x9SXLURZMMfaL7y3kfOgSILZRaQWckcoqxCBygJX/7wOZKjekXiyfe6Zsd
gsHG9tuPQ4yX75NA2WGsZeLiuaYJAIktnIrM5Vl7vWpn31EfTmLoQfo9/sRtF6Fwhd4EkpAjjEos
cAiwlSVsU2x+NFJqvtocrDlXeIyFGigzuj2i6ME/6QgiKN+TWdtONkOT967b0IcC20WJY1HWEdNq
8NnhyK87NedFtZ1i19/1aW7dpplNQItEBIO3aTyAM171UiAICGkmkghedzuasl4dHueWP35EPkp8
JvbP72/SrbtGBFk6Kuw2PkYBnybvz3CcSozLJratf9rnHa6svjlmcN55QI4aLTUTEQv2VzpdgcJ6
W6NnojvWlfbOmXSUNUHrc2Vp5EElKi3QD+K5gL05ZBtHhno0gHlhuMH9A2mow2tb7xNA+HnbSAVl
aSqJ8FkjyEgydkTwQU66UK+cj3tKSA0vtQevifAqYTZEH8icgM6MpbAMKg1q7V/7rmZetClp49Av
z78L8idgvSjBJmXk/XNfkNAZkbmqZa77epVdqNkLE8S2hZgUlBRueUio3fyhIErcI1mFUgoRyWg4
orna7MEjTSalKJYN45cSgUcjkeD6CarfPS9RCBSRjE4NxPfFDIDFRsHO0tXViODSKvlmUOrCveyr
QGCrw3o8c0ESbnrO4cIqSp3RDYHlCiHdEsMh1Go3ZsuROxjjRiRGbrjaoCMrHsVXxIiaG2Xy+yT5
sLDO3AbetlD7t4ko5iiAxNBumri5GqaiuVkJw7LCXI7bYL1kHRHfzIxHbNCrMd6/9kQCnv+XaIWb
FnHbwCCNYthSdbuxDs6z01bkQUKNpi2l3cKfa2gxuH4B5DiZZHNX3Gy012mPR8jLU6DaOzsBzIAg
s/BJ0TWZ3RF4FvWPduLpnuXU/UUsXb0FPyJ6o2V3u6Ouq1/IbUm1pU5HxXhWr0RIyKPz0Vu+Tm45
lv19CjZEOIG8bWIjgcDtzQt06QFcSiI8FHzGYvzjvHC4EaIRbNRsRuHHuyj8oImAVY6GLT1dfov3
eNrFQyzcM6f8TVyRT11Iyq6Gf+EtuY7HfRm2ESTEKHAz51gOtg0jU0do/3rn9sQ3bZdkdNxzsxzs
+WLK+mAixyGbakh6yJbS0S28g7I3GihLXELSPLeIAX3C499tPKncF74Dvx5FkSmnTjL5TFGZ+dvr
ViWUEB5BEhdiMTPI7gHZsNtZ5sZ8aoh7+Pn7YAQM2q/NdWNv0vx+TRjI9QlBhGhnzzBQX6QkOtQ4
5ZTmugF/105Ne56twBVf/FD0PXXiXhdi9n30cbFzA597eDohRkYbhhAP+bxjDplUJ0DFq1rkcK+M
vm/EugqRXm75H2kpV6ieFBgYxRKD9CKVTmGiILx+QwH4NRFn9JzWL3w1/MRGbJuh5sf961lMDeQn
q9ztoiJZ0Sf4pd+5yAPyb823JbVw1c5x41KVOxfV1z+eMvsACb3WaP9fe35ftCIc3uPgfZWWkqB0
oHTkea/369dawt49EDcthJtXqFo+09glBF5hlS8HjaPpwsNOaZMCi5PplsgLIYfidAMOlCVvJJhR
V3t2VQWQcm8hAWfgcQ0ECRiVpt5Zq++unMKUHeKkGcv0xOuvZ0A7mNTq+nB5S6R2Q3C0yeheiyqt
ODpw8pVQUucwWXK+6n0BaOyC7QrewtvN93Lb3zfAr2+xUTZPht1l3qtL2y/Gov26GSqvWRvJt8f4
duZQ3PdoP2SCNbwOLESFvqDuOQc/lG0h2Ot+2qelFQFohaEaizeLGVOmSnq+2UeJihtoTYUZShbu
QMNAdYRBG0kdBnEDTYPI5rZMLH9OrBnTemfj2CaPZA/WT0P4YnU0tTbtd8sl5z7LAefjNJNinK43
RvVrWr2q9Gk3/VJmJ3O78fJ800/nzp5R21JuupNuu6GFPWB5BLs/dw+kFQDvXd2IYYITHQjjwvjM
LgA1beenWcdzCl+09xJseD788q9NrnsNJ1mn1BpBQy94FzgnbfhwSYOsznVTpESk9RPndo+qaPGY
eStKbEsS7HHRhCNaRhlhwoD16ExXQFcnx2ReqU2PSSxsif2Zh6014+mW2vmSZXm6jQSuJ0KMErfr
vyOIS3LCW5o3LRrQhLriSTeIm3N+ngFI8mB5FdUwBmHBbLgGAGS1J79JOKE10PAJw8c9NhTo73XL
NWQ1jinoXtYhDYPivzswvBSO6eiMtcT4a7L0H3d3J6OlcYVDGzi4PUc9LC9PMo/ykMs3XyrpC3Ix
nubOE2EwHq7t2DnOF5KQbVHj5eqbT2Z33dFc+Cz6Q6o5R8NYE+vz71c6OEat0b+C1YshIkqRmnpg
CeZzFOPv/rKKl3bQlaf+I1maD9zlH2CwErIIQb815paEkGs+LafhI3kCVBkzQppmN9MdwBmWoZnm
aMxCb3PIMKbSlS2KjtWMsFxASjU0mM8SLTDLqhc7fpMKgxC4u42CgcNP9gyP3Ljr4TwzX1vhiqYx
r7x/0b+8wRxuX/Pi3r2tE4ZVLQALzx2KKKls1ceDyOwbeKStffddYGWcibgUGcxDSkRFX3XjXU7c
rTjr/M0xMAQMjle8GAbfcNxfTuxh2/hc+2EGFFy4dwPwsLNRWx6z8uEgf8zQUcpcCktxOqbXlOVF
IQPvy7W9YZdYT2O4azI40Mdmk2ARCBAUyJqe8UT1IMY6HoPHs/MZnQr8E6At3MQr9fd3n9K7MH3c
hlTA0PyeXxHioXwFYZCjGY61xJrP581a3tzWCtJwi9R5qBYNAS8+C0AJoe+ywZWzZR6XsWbWKE/s
JfaMV/MEoSXsuY+1hD8qjfWJVAMpZ/+ivj0qcJA5uAQAITUKeat9B8Gb312GZCVXDudz9yaTkAvV
Ywl20ud/Lai3tqr9mg0t/baSfIdL3H1+CcHVUyVGhUStHNakdqhjfDgovVII4ybpmH2Xty110qQe
NozA6bTjNYf4xM9MjkPW0qZ3fRZ4HGVqWPtYm4Q/pcrSC/HDWzfG7zggEMUCx0DLgEUYcAlZhBSY
39dAbfmHWs1ypVaWgBkfyrQmGO+GyyLpB2CER39JK5KjIkXHtRHSsvBn8E4OipMd60lvja7+Mqkz
l0UPdw/JWetvA+E7nF9kdY6OxVr2mRaQMTq+I+9NSLnKARAhlsZmUjwCgT+xpUm4/9FHivI9u18g
V+PUD1z/U9NVi+EeKvVFUB5gNwYMXM7ZQ5PTRI3uP0iIIAb9WDRdKjPXaD/W12v+8kyGUuamWqio
Ugo/mvd+oMHx7kKIYgEB1buPhrsxj/HTQPMYTy4OKWVUtmXbLECSfRmy9DZXKP2Wf8u9YzbM5l4O
LJ0F5nmx/Ph+n1nKarlX19avvz5Dqkjs9Z3Dm0UxQCXnXbbcyt5l3+EYvTmgI+gy3xi1CwSIrFCB
cT7miMjuF+oiGo+94i7ahompbBJ3mjJAwVGq+rMGs4M81uvd3Vc6IvrNDf+wWp/D0xrufxdPPb4O
usImxLO2CJz4KXJB9CQyzldY9Kh54NG5vlZ169atQpqA9dig72Eyv5rjQFbzWEXHClUBe2ZzI2K3
aE4UNpUMxYWZTys9b3EcYtWz19tjjRXY+pgt2YDXgrPItoBqOn4kynWnRgCQBUoFdJOdpCLt3Xk7
THNTnFlydGiZ7kfWmIbNlDjNYAgc8hWXvQFL70wfmrBWmNM/2wv8lmPgJBHjWGfqSJaBzGISg31S
kjLu/yRcr2tY2d16L1naOTpn7hL+bQy1zaU3cl6/CyB1cujS/0YcczOSjcw50PwmcCEMZXpTnALd
nm+f1Dg4lC15rz7J2pA9UQMRDa214k1Xkaahmxe87yGwHbzQewJMiC/a45xYoTvaG3Ioid8EYLZQ
ZRd0G4CCUPMhvZ9flU5edshQOIm8B1R586gHIubmEiPOZSRTbwl7GfNd6JcSNe06Azmy1yuItmRw
wDWgDGykDFkkg47hRgFggerFSos2+pl25L0Hb6BUEamj0q0VGz5uUfj9JruspJeEskNSADm/uGFa
xmYUudUWnoH4MiblbrAMFCFoqMtxWKOkE86q988Hd0d3ZfT2e4lCk6UlZ4L+lLMjJeYdQH/QGXnu
SUECFgYzjtOqgPlElvak8nx72J3vtDU4Qn4YK92tZuwfRFTekNh6+sWO0v+kNH6wCz70RVFU1ClD
8OS32N1wlSxkR9as4oRdLDSLMvJJeeSiQWZ3HHHO4zcq+McQwrWKO9Xbfqe77DlzoYBkQhLRabbv
y77au05lk0/WrrpOJ7P/5auTnKiQg1VfGU7pLk1sw1TNnK+o9lhQV32riDBm+4MrF+HWwnhcs6a/
BaAiF2bfaTNEt5N/ANyifqn0dAhISTCEumABrCzElsFKSnWmgpCng1j+GNbZ0I3NhT2kOcH21URu
qHTFU7gHifqwjDEBggElhTu1JgKn5VruehqkwMmKVkQ+/hn7fBueMB6NmJPwPVC4BgXRMW/5Qujs
UI1K3Uw9z2WFnfW9T9JETy3D/FhZzMaugcHe0uSme9eUJWS/Qlq5iIT91giz00UfQiuCl2KcnA07
pfxL5yKio/zsB5elx672r8iXxY+5E+e4VLVkEye6WNC8u+nooFvElrq6TXQbYwq+lPg/K9/SsXcG
RFrK7TTBxQx1SwLryDlaCJlAF85TN6HY6DiqNV1uiKf4EiQq251MmMlLcaG+9+vWwnXEm0sFNoI8
FceHVa9HIfyHhdS6BQZj1XR4IuT6sKFwZEqKYkF0bnpqbWegJTQhAbnAGjzNHinDtfY4XiB8SJHX
jYi4KUKPDu28aSlXc8mu8fW8+FfMnWR179LJE0YEyMreaB8Nq6Np8cnN7qnziE+ehJ6OsyqcqIZ8
k3s1h/pKngbtKFuerYDdyjYmnIJ2t0KIcSWynqFvzZP4GxX2yP5IB2zo1Uol0vgMLNGBFXHT6ujz
sxRmLEdVU2zbgbi/2Maau6V3cA8jVDOTh0FN9zSzJ1sRbzb2lhb2rHxepqq2J24YvcEuSNrlBpiq
38DLnvu28qOuFTqtx8TrUmTIKe/ESNOOp8qIDmwyAZ/fXHMQVpMRMSecw715o3QFxhMgSS+aLF42
cbKsWlull6SDq9jtm/Ft+xREnyxpuH7n9ZUVNqEbQdCKXng+CUO5Dql+rXgayCb8w+wVMb9RCuM2
pQIsC1aSzOdTsFPqYHjMEvOOukouOKgq28fwewVZ//BtEt9GqpuNGrbjn+p0XkKdyXFsoaGGSa4g
FH8i4AEgxz/Lbfw3auxhQjfPM7Se01UrUFON6vcViOw3/I3GcDcVWaXK+elMr0hcmZG/obhWYLhC
KaagZkW1nT8Og8BxOBocVFFL6z/BL/oQ9ftbb7gifnxBQWRZLZh2QaEIl4IsjC6D853rmNKpJ7Ja
jRS08xRG9YlJRH6mVKgZhJfJcs+BUeKdw/RJv3tWT7suJ6bdmy1xkNDQF8l0AEmDS3sIE6VznJHO
GON25zSJcIqzfyVzggp6I4TVP65xBA5qPgY5MsjVcoU264tvdSXl+jBvce0lGN9FKXXp1QFR80yE
5gy35NpsZuYLGmLKdBakFvVKsyNX3oGwPCccuVi82mMtzX6YFAgkEe/lflINR5dgaWOcjxxzenl6
KcXdfBxeQPODvMey16oG/GRhieo7aCL9d0lI+a71Pa109Sge1KWxtp/v+i+N6JjS2IuKIP73kJg+
3PnwqzTRt3yQVxeQfQKA0CSfvI187DPV/fuHva3wVFELAabDs/tucPT0SfUVD5jAAlkJHxuvC+bx
BiW4ew361j5ynBKEC3QbU09UV89vNQO4J7hSA3cjcLG7Opn4rK2hoeFYzv++993MlmkzoRjXdnKs
t38cxFPX4WgIbKpedd0mJ+isn//Dq2qYPNDZXzmCJS1f7NSnFBAoIOk0NWMgX0I+TPHVWOqvgeXF
TE3+lTefQ2W6LeBkeTrNIuz3Gl2isBSZ5qIcxJ1xUUBuVOlqL1gZwlqiaxFo9hD5xVzzfRPHeT5+
SUTv0uLgyxAUcM8NI1dTrufN8fecndmXj8mV1Y2Nij/PTa+T3K4EKbl6L21q62DRg2li5xCy5aJ6
mH+hChZLItm6GASYF2UglJbQ9ydaAClR9cjHn5KUjdXhoa1DaibXDfuyuT/sV5uaD/zUncJ+URnV
kGVaLSyJvMhKx5lLFdCxZGcXpzrtNGMziyCiQb3Xj6NiepJayw3HDxL7jOFLVZmTuMY1pL2JxFOi
jFtjedok2AERC/k2IMN1Z9yPU8Mu3f5hpbH7fCiWtAUujafC8PPZM7MKF/8a/7p/QSHNqRNkCj0A
xdmhEMybgL2VwntLPPbfqLdGURNbNMcH0BG0SCPia580aCh1bMylmCAWnFAyZs6thNoehlJ+3Gi7
M6L59LUellNecoNISZq7GDlg13jcAcUcWLBaj/+SJbE40G3e1RbNQAKNUy23u5HOVPlkvQEyLdQ2
u5QVnQRnRTxm9U76y5GZnyLMmkhvoG2yN694WUSNyUXB3ZEfq2HkABs0w3fS3XeE4rPpN+EQ6Fis
rNU2XaqLkQP7jBVeALjHKKYPc1xhhjQOBGOdn+JN65q1qfCjCpc1F5DaT+Ri3ycB+//3WVPmXOr2
5ilMAmhG8P68P2rgjXtQ+/NXcWC4G9lbcj6NPn2ZUFAw7O7dbOARF6YOAwiatB0vmECluGWOgd5R
sdpNesuQQ4UiYBKUxBDsfsxuqswzYuDjJLxUZfUc3SMMTlHKNfWxHsB/pmQB+ngAW0Hg7o1Ocj/z
GeH7NQOKUQ83KX8yGwlqzL1Vf7SPN1r1tp44o80GTSAn5+N8Re++vo/f6N9Z2/7mPrt/fs/SpVAY
kk04V8/Aqv2m6ErW+Hj2FphgZWc8siOQ1wCiwGTevmmciUTWto+777cwhbmXezw9NwHP3/V6hl1e
Mkea9dhPKZVXpvKFgh3bnbIv7FZbHN99STK8DUqtunDL7CqcrL4hTiJ4185ouLhEy/wK/37mPEZl
kHKDNFdxH2lGxgrPIbfMjegDi1MV0OSfrXyvROR/39D69i2sVl6LbRhtCcJtiL4vTq8Y6eQYhIW6
bQkRJx4egG9fQG6EwaGkbYG92++ilrB5BVunX0GlNGegEuT7FJ+rJtt9V+eGEmdIJkY2FziXF2B1
15kuEZKWM2bJ/7rgOWPrWM845Aqnri+gErqrbh5UpNCjKOiEn59eLgt/2jxGgJNbUDlNeKr9YCvG
OAA2F7yh6cB2qD2BbUU+fAcLQZ2qxveZkV5mUETIR+o9NKcHPdakO0/pNMv/Q9EJrcpwXq9n2HrO
495QqsxYOQ3EakpD0vxM6fjeFhRP6b9XORrEJy06S8X60gTiOujcZR4/iOyRtDlLrHT+YqW7YhrM
9cbCqPrdCowZomK6pueRHa4Y2ikIav2N0aMY1izPYZ8fGIprlDb/k1uWdfbMss/dcbEoo446e7Ik
xB46L0i+LVPWCmrPmnRcUZeJICXo2QA21GQ/ONaq/j7lRTozP5xO0oKHFtGba9nbYa50d6U2pUjv
NE841b+N1ddcjDmEZz6Ch5c8+11Ocb7V0RArEGd7SU8bTxQZf3HjZTNd2fvOP6dNXQb5ttz92Q1z
z45tGPFEE0l35RoudjJ2bqJCefCfCJ8wcp4HP/0WtZIMzO4+EYdF0OPreOIBzzyNUitws65MT5ZG
zk+HgkT4n8SI7l9JOkAzBTMHuD9XtkB/q1w1Wm5iL1orj8wHEKVA0h9eWUdZSsdeJiFPl565KkGU
Uwv1H4ELngWzltnBVekua0pgvhXpyr6Y9yncMpMArGosCme76RoQ7eR/CnocCl0E8cUbmO7sI0Mk
KJmAa+Dd92bp9gbajgcsnBCLkNuZVnonoYSEaQ9efoWKrrQHZtau/SZMVBpZtVbmXkpCMumTjixc
liowfo3zrvTD4ZIKDebtlktWZ+Pc8zlyFsI8ux/GGabrODrsTzPN3OEkZ/6H05sU0E8NQuDAQJdR
BekNspMPP4Uq6YwGgRtBp1SlDKdvfXBKhcjdkxkrbviaw5q+RzMR6b66qvW+JE73TaAvdKVuXs2b
uLgAKg7SoqV2onqOcxetFA5m5MN+it60YTTaldi2otoOxE0V2IH7Qc1oR4b9MTyekgR9vevu0qEi
rarC/NvGnnmBAjI8f+zwpbu3SfLJ/ERyEJNJINX4pwUuy92C5XU92YHjBRIs4MqIJMYYKLGQVxPP
t/H4nmjYwnOQ0UM8KYJ/qz7VBkI7WXMI+zlcYUbAriK8850QuiCu6oz58kwN1yn2Y9bugubSTKcA
AUIFAA1N8nKgwH1mQo7dqYKC9sOVlJ/TzsYAyziJ9NVnM5vSquniat1TJCrVuZnYdQ3P/5Q1Avr4
q3M3UEA6mejA5dTGGLu9W6jnWqka1I0ychcjVj2YCQ80h1cJ8K85fXvH4w3hLQjwvoi+di1A+Xrb
31xc3f6INFPIxUn7LGy3XOfWyPV1dGAuYmB9uqm50nozldRBcQS1xjz9XNWAY0+cclCoNqNZjXtw
l3+fWymGJ3G/pQ7QDjNwd5gunriWwWZkNgTaVOAuz+R9B91qDI4BFXapHuPy8RP1pyVYz5doEXk0
imBK7Difl7gRE+pGnTkUGU7/dwho1fJwsqmhEaceAteznUndAX8AJgqyQ96tjhrCdmX9MA4ZP3qF
6O+AnRHI1WhgYsMgGZDDkygbWpbsOC2LWEL9SUSxXJyLDIgjOOoSHkRIEHsAn9sZQfdwwpf8En7b
1M5nbZ7cQ8HjKiNTTmjAsP1Ys4d825J01VU2G0gNPP6NUjHpazvGgno3B3D91qtPnAiL052X7kFd
HXdgvWqa2yygbmQRJOo41ED03lvVvPsQ2XfbDhTZSWaQsfnPjq7YHH3cV0sny+IYr7Z5sBN3ADK1
ksueUpGb56epOdaJIPkIRc8dzLZUGI/pAJkuhY9CiDKhrBFEFBq8AFljmehNNPZiIOHzoVNllLQY
bkGYDTXaLOhuX5YscVaKFSPsdYOXT9r8JUPwTyk5+ANUII4c7kbwIK3eeP7z9k4zfjWs/vyscqrZ
TLED4f0/UXFzKtGUuFd5kFUBl4swblVjOAfFNRuOnfTw8pGUWufzOLXH6dFpzRYDhiiPF+7HVYui
/XTHOSLAZv6XWW978HhP3+qxC9x6V0oSvWcYVLs6EhnOv0G7kL+/M9oqx3M6rAh+RJf/zTNWinnB
G+HKPKDqXacS7jBVev8Ucs+SFu4Av6K+Z06l62mMsw1afFPlBG3HYajobnrX/yI26BUYtrmQ2MpF
K4FechGjciA3Leka0wKGcvVgA0WmjoW8UYQLQ94wtj2OL0uE8c8IFjt6IxiBbhiXWlOEul/+kimT
z6GXur17+F1b37rP+0MsqUtLMWXr13/Vg0jGi20ZN0XaZ0ihO6G3tHoI0I3tflSk9e7XXXyD3L50
AJZtG5Er6kaDGJwqf2WbK8Nka/kIpmdIqNz/BgXSwJJdWaoUG4MWLHJj/W0IgFvqVxTKuVKIiTNc
ICWGEykbRQNfHjmVjY5sz7b4yfkfQqZMzM+5ALH8xNYoor8Gx2OuPOnFxqDzTPk+fG+Z9uSy4IxR
umTwXjIc/DuBlEQvhMLPj3tlN07sKjiuDtjXXOqwXOoJFDsaPAxaR5JN2Oaom3OrbKEnATm5wROH
IOrXZQDPkuZgSUpVk9pcRiF01tStxm1uwSysNHiYBciAY8ueC0FRs7CpcfYAnLXRIuYpaPmm/luE
av7SNTtR/92O/rCQPlUwHnXe84DB5Tv5+OYEOW/SqRmNuDzSkYHg3ouUSz/rh8EG1/4Rn39HIrpj
loqnVRGcGDnt+m/vZH/U9MEZRO5DO4Qq+P/S2y1mgEKw0/ZnpMAF+uxIbVUp6RoDhjS1Kns8ZxWd
7tpTMhdxu51FVumefi54Yuif0kXuh/uGA2qrV0onmn29Oh76tkglcgdZoVDqktzQscyIV7Qo//jG
oDwAPqSMar4k08Oy7pa0+GWBZCrrRY41KZu5bq+V1Wv1Zn9qrnv8IfsAytr0tuTddLaLJM0dykCS
BwtS/M7/46FPfaGQjJCLLav3TzsaywDHJ5iMCqDiKTER1N8hVsVO2b5pn0sBZhYhiKCkRyEkByeJ
bJNfRQhGl/s3/jR19khi59/94nw6YqNtEzlFQyXovQC23mSZ0thH4vNfvpn+OZBhayQvX8oiKQYA
9SVCKlHM7oklztW0iX5FkeXmChOFJwUuxf9XNiWA4xrF3gO4GWMrkccL1ORLoJisYwShZv9GebHc
dmqaPz2kJ88i4jECUUVhv33IY/4U7ted8CShlsHB1c12Bj/CcUZbcbSd5xNtNGN4IC3GgF5LxHji
+Rai4bhDOMSn8VxW4J/bo0NiIf8nnSdsr0zrlplZKI0PN6qY9x3F2YjrnZ9vpx53nK+wBi5P6wFo
4IW/HxMWTX6InM537bFr1jkU0K+2Gxx3pDgpXCOaOh6GYcz0Webvh12hsXuf0Xb0qz7xXfM7cPZX
DiZ5mM/PxcKqOyh4GLwBxE6hsChBNMCVxGahChXd446VD4V1BTOUUJvDfUS1BOU9R870zL4SwVzE
9TBEGVzJOmXo4AmPBl8kqrm2z+0kXqPuofbzJRXKBMzU/6Ld/gz7jxgKz9xOw5UjBSJ/ySAK2c1x
E9vQx9sY/DAi7FUOr25nlxEtyojC8FunhZ2h7eembcJBLfRRlM9w6//kBbcAyHijK1QoIACUKvOr
VwOVDnPPStE0BI0zZw8nk9RKJP5M5Q4wv2T/GPLgVU1/k2FwweFEFPWuDMT54LOwrLolVrnzG//9
hlvVnJZl8l1T03jouVcp2MWTDTIhuVJhoN9KlYUn0p8ASjPPLcxHm3ZTae1NQogBzCR9un2hiXhw
NdhR8pFci7bly198TSo2zSd+LQnw4ercxdkFcQsoXrAKeIlrt1GtF3CERwN5Wehkrqhs4KTjYDWr
fWJF67ny1fiiyT2wTtkK6CULSnSMR9Efd6JEBJBAc6ZVgGXx9Z0Jj5DZa4/6suJW2fm/D1sPmmaM
0/Ex0wBEFfSFspWRgV8bUtK+LG5Q4bBN26Huq6q43G3w1+UG3IK6StUGYGT6VbknbgtkcBCjqaqe
HD8PZvTWLtp1o1U+I/dHiIosdLJnZkVDRD9KRphTYTSlQ6KHvZVF5+0vkKRuUDdfOaVuBBmpUinj
PgCoLSF1eMJ6ENPd2AQbdjnHXGkwKxA6ffwtXohawHfXwZBnzBpwAh6Kx74xP7nU15Zs7+ymYQDO
XovioFNUqlsljGUd2LWQQcfMeodEYVKQdABX938bj2HTaeBdSgw1Q1fmcIw65FqQG7vrt16eTiOF
45LhJh8fwh8HHtUzEzj2W8z3vrLZo76ueUmkY6SvLL6PXMh3bzIHDVIJnU8r9PWjVh6bR65yTWiv
7nK6FJrEaSjN2oyxz2RfVLwUTCUbHhHo3b3Enjn7v4W5ZB4xiyhIn0LPEI6Oj9pcV3yjG2J0GC+a
O5qIlg9yTKdV1v2rXKV8TNFsIRuoi678CsfQ6K/KMGJcVfCLmYesLEIrYbFB94rETVl8R1lh63KF
PU/ZthqZ/BN0u3xeTfjl8/J4L1WfVUkN09I75ekct/tjO/75A8tS0WRFzJ+BAPq9isn+5iPuZqlz
9GpR2DUM8c3+Q+WEbudPw3sZYoSovYyawnKxJooGrfwa6IIGQWc6oVo9rNZx41ldB47GQEvgPKby
VMkELVlOXLONLhOxTLnb8FCcszjMfWJDE20SxOZUU+edxtgvjNXbV1+0t7msmrLbOBzXtPdxHcd8
rQLlWlQSV7WjimCgZJXx1QfiIkpkLZKCodfPWOTQqWyprPLJ7+YsngYIg1KH+v9huDp/Sc2R/b+G
DCkO+/zGAj/qyRw8kZmEH5jNRXdF78KOhoT26WiC49m+Wn6R3WdOCsZPOuR7W5iEvZHStdwuJjK6
YAPTSpFXMB9/r8o4FpGsEdeEcYmNmeD1CZa7JvOpwJ0nYKAa24m0UeUmIbxm3XllJY/nduofc53C
PYH7SE4aGaDvWoaLaqp62TQkytNMw3SgiwHufyU1yKKI6n7ev6uZM5SGrpZT9XXJWmCYPdM9Lf1w
90cj9X+WSEXQ/wjmaES3h9wn/6k58NaBMqUfpbAZimWHWcmMK2/JflrhzLpen9JU4XKajkYMqwT3
36lGpPVVA2x/2wEe7zkVCuZnR2iz81qYtQDyVOuYGV8OHhWd7nFDbQcfEToyE894TO8Cy4jF1Ayt
QWoApMuQ9XMPHYAOR8m2r8GYRvovV9PkcwwzFYkp+XFl1HklAGBi77IbVRMYYJAA1bkj8DJxzNJu
RFvvxDyO5pTy4/YWHH3YJNpr0cfXs5HObilUfTOHkYUaGxOVD8Ex7sByhCyWEwSIeMLgp4xT6P3+
T38+TIcar+VgS7U7IJ+GXdlOk2TYXJV8rm/gKD/0W4crW4SDceQf1pcXmtjJ7HrVN6ZRy8j8k4me
kQyRiXEAUf6dDFKjwAKB6fwftec8mLLR2JbaDE/3agLa96WpA/zcfc5L0PtSJTm0H/8o3xDFv1PH
CpIDH/qwUsib3UsiihA3q8A9CZxfKflWp2uUfhMmKPv3jhi/gqJbm65utOz0kkkafFch3BNRbTLo
WJIyUvvBQTCWFBWz0K23phH6Vaj0ckGojL4ZaU7aC8VLTQo8+sXfL9Gz5WjpOOrA6fMlwdGMm+7+
bpyofFxhXhiKOf3EJWrt3zDjS9LeQvcgL4HcK83Vg0HY9kSnq7fa89GA13pqEyY6833oC4BJlMCX
s9HIuGNFB2PIEm1haPwjQlz9yL4YxFiNQzNGxmgcuo7piVRXVIeJI5dXpDKvI83tc5Mmn4rSwOVR
knm3qroi8k4BTDPSDnLE3KUE02NUkN45h00RTpiC7hSzE8k3n7gBMxguHVbS3vuKFnnF5JTpIEaA
tu3rhhhv5HnMh9SuhD+gy+o1daaH07b3QZedf9EisYQBRzGtQc9Is0CUyht/IbDs+O3Od5Mz0yuY
I4yBdOyFvdI9Ttl0d3OPpwt1BGBvTBhGBlN7J5B5PfCBekfurVa/bVLS7qgeoT41CAVf+uhfddng
SlAeRxa1wvyU2kRFWqIIcUvCTPmU8xFWTJBslQrE5VQNIUxp85lq/6WkyAVf/KhwklXXDe1QWnvd
L2GVuLn1m0qpxoJJiIXMXIE0OlDk7jj1pXuQCGuUYru4IuQ1vAo6L6VCfXy42/OdKJb080PwH1ES
PBRUm9nBmQ1hvZ/6WJcyoYrEjEoNz+A3AaN2JQTRZiwV+Or5uhbHpxe5s0OyfdM4lzKHa5m0B2AW
GHsxzPr+jpQRGzKYk9e7jds+CVlx5kVG/tgz/VTJQdkCYXa0DEOgZFbiCQVf+r2lI6VoYzct+jxK
xQwarCy3NZ355d2nIZPTUZfF4ojhJ22iGNEM/gnkXl2WU2MmimZBVREwDrxHG/MtwHVW8W9mKxR8
Wocv8X8ne9Ssy0xPSxSVYivB0vEKnJ/STBXsKIr5nu9/yLsq0pXeQT8ZH55PVeik9L+KAeoavHhh
W43qrc5FVs9olKtaI9DIT7TJJJHs4gIlcWTsM57trPzPXpSEF0YmxqwTJA94OEDsOzYVS/6pkv6C
jD+vNUQX7dHcehUNl4oj+YetCmq/p6elNwisoz+tqIIQPzBt+AcWTZ90Uf9O1aURgWi0riKZjbTw
SlvKUcJyTajyQxAwXup25MSgdgkbBzt2WdYECnBvWb6+uWsIff+1EGgsBG1nIT2vOWFHetnLSxJJ
PfjkZZsHV6a0ZuNRU8zxUXmTzvbsMhAib5ezLhEJ5FiXrhs25vDLjQie9eZtaZWcr1AZ8tSRaDug
nPSPKrGsy537ZSvaSndxijiK7nwTLKh9XQm7APVLhLYvWDstZHWWkBV31mJKOxTpR+nYqdVzRyCW
ccbT3nK7C72L0STlQcUov/y+5ibdmG6GDWER8UFajKT/tHznH6ElqVZgV4i7uiRGm07q9eDOGsm3
K5bssK2jXdMk3HOrGQ9yS9ciiQF9fMyLOoubvcYf/TQCLX3VPY4VTxpL48Deozm3yeHsB16pqj4e
TUkoXEVlQbGQiW/kylJE2m+e7tGumMTbcNSbti/a2z7uefOMgbHSpKgibi+XA0+Ik6/wtIh4ATKj
nS7uRSsUPG+Mpkw/xmZPJcQV/MOAQNDO2NEr33Yo8K4JALfkXmT9RV4/ZOTYtQvaPnhtt+ppE2Ea
u0Q6nBAzO3ncH709Qni1sJgEDha0RyU9IkYr+CwgP4b30DhE6a0U678J4GkEX7Qef/6lhM553dOG
K6Q0u3ceAY+0dvaoHd954JQxSC19yjmWONtCXCGIQpHVtRdJ7C+7e4+kZwL6gpqPe6M1IfXPVAUz
y5S27TEx/HRSy92duzm8Xv6GypfghXWRjfqwT0vsQsuaxhyK3c0ZcnRtEHbydr9YAeW8wcSKzJ4n
nH8gtQRwu2/4QJGteaiEaCltof5MhvszFVdGzTz7iBAjPjj347cjc3CCaDNht22LQp19lptaYjVg
vpuNYPMhZsDUeGaLQnPiXUjLQ2OMei7z212qLo8SIXjfLfwikp3gDvc1eOErCaiC+lIAeGSuneeb
CeltfoumYY2r+ZGSd6BEF5CTHb3FK8wEXcNt6ZwG2CLrUJgr2PA3c5UsQZPuR68UjGOzwPKHYTLY
D280oC1mxVuK+Gj/U+FrDAdqa2GL8Pyop0Tc0MXxs8w65RUIX7oFrulwokQDO65QjCJOCUNPi7uY
rUrhglJaaHKIj529Tgkuk6XBaJtRshM6P+xrpobY9mxcj3so4lNzMfO+yTXTAHT/lYWtoSgA1VyR
WoRxlGOSlxlm5VgXri3gcXmy1zcW4TnJkHVaL/dZ4QVmzCCLHvUn+D4Pzo30uiyvJ2uLzV5SPboD
30hpK2/opsdfbFTjv4NwQGNItMI5AKxyrWvZpAr9zKOZLBgW7PktXjrBJeOUSzrtAOL0vLhAsmC+
bVLuHFKMNgx600/5oD46WATsAhRWeIacXcD/doRe11uPfwHU9OHi69Dejd6rQZAqWRK3hBk+1dz4
21T1IgcH0wO7WyieI29sKsd445npD5cE+QeJC+f+AjrV3hDjgePPyh+/+2cHe/HArTt2d3SVUVLI
dTGw8pBbPx3W32PYvnKnYQrHV5gfTnnbKbbB2bAHQ0RvXcQpkM37Tv1uQYTlttA0pt8E7io83ngW
ys1OuDjVuQEN4zuXtKJ79T8g/VS1GMogxJa8S21g7zXQOg1XDwaDo1ja47/koXPUQFtgV8FrGVhi
3IWQfBkAiAoJPMM59ZgFi/dUEFQb+Mc5ersus+OhDsrEGCM8l6xYKc/zDxLgw4/mRdx822o6rZlR
ijYBkmOxcXJIHcvNUub7qWJpElkpYTAmMRSsSNB9/MfuNsOrXMZGi03j29I1ZyuWlrBOqhkWUa5P
ZZRbwCH3wX7nWalKElL9BQ+IN78K9kywWNGtZyU5B9/R2AlKideBF3NO8tQszj84ge7uMg//eDQu
1pILD6hGiIOmq3uCWMxnSnwd8VODFE6KpJenMgX+fpoBuYPaSyQWSGnHsVM7Usip6kvuzmzeX6gN
VJ7I8IQQkn0CManCAH/whlKZKvSmURmSIkDj2nsZJq6NuTGTWv74nTwwu/Zo0MpkXlUlaXePeBw+
dwdTB7GNTsMk5KHvEgJ+Fxn9tlTvf0pOf1wmQjSqJyd6GSdfsWhlDPIFd1LhhKLJ41ygjd4FDQGc
z0uymWiZUnOmm8VBaWzAbOXrJYtpYR775qLE8GbU+T/eDioC4Qi0kTXZvh8JV/Qyb/SZWuiFe7qk
OFjfozzFYDnOz5o96weOq7dfb73KJYWjlQW7Q3zjWneLiP4gbfbkAuj39OmplhHoenHsvWJ7DnuF
Bm8svReLUDm1MxLOERMRKL6/213hND1BpfkSwOaxcON85NkOEM72yxS9axhszVYBZkXBm6JM963n
XlV0gBpVXGBFnLe472NuoH2CsEqxij9uAFZiNUJ/1zxuaKjRIyhS1DNBpFT7aBDyG9DpcjMkCMO9
4+XRVtNwJu4M3go3I0CQ7YGscXryROjGMOpZoaakW4DHrFyERZqDujxgsSC8HKkIrxA6naByL1b5
nNo6fgH5jZekRnSGlbbCf/EwbhF8Wg6fw5Ip+mi3jd1h9asqeoJq5qjj5r6t8k2tMtgEdjGGD162
A2okGqsco6s7TGGjCGl76oMe9knpwmiX3FPJEoIiClBjq1dyvZn9cosf9ZK128JvakbwwPOwx+Dj
LNH9vhhsU5rS+ew2t6zcB+o+DCyKkrGjDZ8tMXkzEBoIblOVlvhhpJ+WgGub0OmyBGMyJiq++lnQ
qJ638qCceAvU402OkhMA3yGkr1f5EvlSqjS9tVeXH6nroUBggwtf8KF2zV5GQpdeA4FKUksx0j2D
4J9i3OtacaDFqwbp+6SPjdFsmDIoKRH4YqVqkJHa9ji3VrShfpuID3Ufh8fP99UrxHJVjuFD4aVs
NnBKZXdfFoXs1ztiRO9buXlnqYMOxEWSAr4D3bL8t9fQyj9OvOzx/9ZxLi2Eyp8x/v1xNpycFo+R
fl74oxebW4iLa1/8qEiUU1BZWJ1B3MDKpyXUKtesLfowBVsN4cZm1mXojWGaNh5vMb7RYU95vjpy
C/VqWj+klgvg69HgapIWXVVAav0/+egUQhetnj1h327n2rbyg4N04uvNM/M6mck7tU7FYhNLC43G
8r8VfdRJ4A7isG3Krs5T4WTOhgjpKhDFz/GYjFiM1acx1FYnvhkVipZStGxKSW2rkqpRS9KpJTds
pA1ZXIarUXieQlAK6E82Owy4DzJV3Ga/p0csEBNVbjj1vkAoemUWFmdfVioL7esiN/QyCsjB7EHE
Vj1TuqE78ZrgD845iYLZZvaNpFPoudnkN1p8Dz9w0xhE8sfUnlSBb9TMhzvvDztBqUex6X7H6pYJ
ntTd8rHUz3yzizicR0BYRisF7ulXb2LuD/y6E42vpS/Z8DDZe0tPTv5GGKJCdPo/dd6ZsksEdaZs
7dHtJnAKfO5pMatlbtgvTZ3oZt09Z21M58vR0RWL/JY6WdIWgCgHw2f3t93SD0ZVJPWwd3/tQkpZ
+rU45CchdKVVzPffPzyo1tLKZtaXBxqus6rLKdZe9jGrFdMDuBVSfSgm0Ws4rM1Uw8G0dOwNGlwg
VRJX2L5RCZf4xhdLci5faejgAjhGa4SBwfU30hlC/PwajfIj22mzS4vV7bEAo8/uWMdTawNmr/yH
vjHVEZXUemh2N8BbqnULdLqM+brYz7Ph1/+GhuGxwYy7aWDmdYdEuaGb+KsR962C/VuywFbc6+AV
rz8rlnRoQoHApZFU02OOt/LZWmhV5An0+9xp+hUDtiY79v2uRyn+E4RS0LaNfinJ4mVzBXTwvGnJ
DgXGVaNf/1kc6fsV41zMJtfTpz4UgocBZ2npQk3KfXuSzCL4k5piW2jyYgqtpjDQj41uWhgBFbG+
kp3HLMv4Qv+yXbPnQSQ7b8w+ycVefGhzDMLEmUtdlL0ex9jfKRih0pdcO/SntNqcOLpF5ny5vkav
Lg1t+9fNL3MXBQB/oxG8U2bbLL/C8YLCH+Qlz42xOmyjlvX/15v+dKoUpN4HbX4Xq7iunpDj02C4
FxKGnScPsoUu+BQUv9I/JvB56OK/Ucao8krhvNtF+FVTR49syKj+XLU/SKi2NsSlujUIF4UPCn/t
faj2QXb7kV8/iVQyuvW4vdU+aTN1OXiWL9bCw0T4aslaXAUfqkmoBijS3lfaGuqkHw/2BA07oy9D
sxib8CYwkAv2d8oB1uTeJezoXebZPKDJFKruQhF0PFlebL9O39GcMVywLmW54K0JZByng7PklnMO
R5rjf9j5ae6Vae+Jf9n4mWuCB71bMHKADP1Jn6j4kxHKWIPObpNn3xmSRXJkc/9a0+zg0RMJYTr9
bH1i0BEKJYzMSkaQy4jcJEQCcNaYfwzNwhb9S1oHRdpRy5C4dOOsE2Tq9Vv051qMc+hidGMFiM0i
X4rZUX1Xute2Kiq8zJJjTO/Tm119PHXgzqIkyroNWwTjrMqi0hsxzjOec3IADE0jFk/T2UcpxlYq
Y5X1Kl1GN4tUr+/mQJLACSHK9whOX3MjUJo+Bx/p0ptQNkxzdLn5c36ft21XgyPW+z8OK22rwtsg
KsNcefW0HZgjO7c26A9sykZEdEl2di0Mk/D/zfVledqua90r9wlG1XeNalZzMgdT3s8fqR0awPdr
dFSqARkVDZe7vQ4NlQ78HCOVQf18Tuw7Jd1wbNNcxsxCsLDXb0jR3HO8p5tRID2OS7tRklafv4Og
wNa4vqFzbMOwGGB4jYNu3sNShAkr7sEW87KlfhAbEZFa4G/umRafnERc4JFnUah9M+YjLHgXpe66
V6eS6WSmmJIJATtSFyzoQ06teeHkRmiXmDRaMyjymG/Tx4BLG8Pz/sR6BHDb9Sq5PHhcGfVioIyV
iRuFeJ6NjbWWXjU/udE+qsdVg7XNygaEuAM2f205RkjjyH+++PUZqzUrqD/p9yTS7FhuMWAF5N0t
6hMFB2J6XXdMMbNaTstXh0RFK5tT32MUO98eUGzgT3N0SyhlOQ+sbbGpOu0Os2Ushma1BBA1mTbW
jVdh4bZgw//2Dx5mUuEPe492B/0zN0A/Tz6JTS9Zc9wSxiEbsn+QW1vY5OarwqsjKVfYB0jjc0bb
0DXWN/rLpl1XCgQBLabnQSxqI05h77FAZ0M2lKMi3cfOr9zDwplS58fB9UDUJ8MdVd8dUlVHJFOG
GKGlEl1lrZS6ZDluxs56J4XaQBBYvEMDHhlenPExrNF9yzWTzAmlSimgrElpEcf00yGjtVMl56cz
kE0C7bvd/N77Cug/y+vRD+aqIAVwPgfVuRf4dd3eCVhhwbeHzr/Dwtkruw3DeAvqKwv49muXRPxH
B6eAWddRqR+QioP4W1J4CThEkVwD8mpu+PdyQnFTx/Z6/dbP6fRe1SCt6TeBA1O6UCkLxucfRfGV
f7ErENrdVG2Yq4mcDlElXXu+a6dz65kSfjyU+lPW/R+48VWqlsjBdDW7HljQLckWRpQ6+gRg/2ru
IShRfKtFBQjbLr1NfbMSkfYIDuhhpe2NRbX1WSDXuodeGDzCLxCKZtk+cE2/aEqyXeyhT3uw+zuO
Zwotqe5ngSpQ2PxxdEUkxb25isyVZ+O7D+aBlQTynnxqk87YQeSUDYLzNBNiSfSkq9KxiXmHg247
3BpSQ6dXys6b+xDmFumm9xtnSU/lhKJjyGAepkIchcU6UIh09ZI0FbTRbwz7yWq4hy3Kj9mqS9RM
u4SgxGztOvGLNC4MwVTCSq1sS2/W+SLLSoj7EWpTv3ur4fUQB161o3+fYNbsUGE3QA5Tg177HU15
ltwOoPr39K/fzIjKOe5G61luc8a2XDLnlE+u4O19J0Empo5TmHajHg9PrmZUb0YlxprWyPFm6Gs3
z/RQzpYnWFjcEEJG7u5V5aeNKDAqso2vS3ORO0/VqwVJfx7FFceJhDb7DTs7YUdPtA9yDCOAZmz6
MVOU4KFFPQT00CuU/ooWbl6AIjEH+jATLFKefPffDSVVN/U1K1t60AUk7OVE6b6yYHIRk8N65c64
SE0FKJgbd3w+M2Y1Tp+5PzmwZRYODoe+CptUfo31ORujQYZLBYhe5VjGhs0kPl7CKwV9r1dYtnIG
8jmdgHqFEsCnXtUftIqp8vzcYxlBWVspAjTAVQbgecOiDUjsCEbAJffGZjPPDh24PNhfWd9mY4fE
uhuMEKgEfAYzpZ/dnB3C47a+3ZwqK5EZooGfBFQY5DDaRCYLEMiPHbAEeqclfwjfKtWEkuFTY/fO
8Z31sTZm1AMZS1NShZqXd+Oz53Kq4gM2YOBMsZMRd46A3pSF4RNT3swSIzxGhCD+BmY4mb05PGA8
HfgJu4bi3KCFm6IVLx6BCiHw9ZApSZqN/yBNznVMJSb2gcJ/CWDxnmi4inSbG/s3V1mUtarvRJJl
YNu/f0cxjW5PyWc4qwqJduaHlZ/n1iCV0lF8BesRIzseeeD8vNRQCHmZgGTHKASvmAejhazeFSRz
gLIqqJaiIwNV0jqHmHpklU6FN3oSdd8p3dC1KiieqoAJQZYu8iF9bkMU1KptGc1FMzkoDuRsAhda
o6AE+JnUyFS4qIK13FL5uVDx+ldYse6K12mayIjRVTYQjSK2xsCni6M6NBniGm4iYwWXTLw/7YAl
5rYa+FC1j28TO2xrSVQtarqKBFOuUot9VwVTNY9PTuKxL+aIeXgN3mlAP/aIk8AqR9BC1IOn8hfY
1+8lKlQbAHrKVvkhwoMdCTLikxLbU1kVFb9SlwTZvDtSXLmQFFcWUdlY8FNHPEtFpXd2ipy5IieL
XafxN2g3kWYXgUl5vLvP8JNUhV7VTOp2MH0GBiMGrA5g1AZ1VBf71C039HmZOc03reYYqNoWQdvH
GnjcypVMsfQO7kI9X2Rgn/t+y/ix9KzCtzb+i+cHgDbUpEJQ54+OcUuxH/nrq6mboJDRSN17kyOS
OF3H39VCpPaMjjl3DwNxvM1QwsuhM75ipeeoGOX1TxCd88M/PwLvxfyywF1VTawGZaFxsdoaGanQ
vSUy/k7v4If0woi4dw+i1Pw680oiuJNgS7kGJYnz2eZqkypImL9/7zxxtPwQ5vJYzR3ltpFWw4a9
F9VIzdQ6DGkXS4blEi/s4DxAqO/taRc7bjBmkhAuzj6Qb4F86RQ9xuAiGb2dOq08+s+VKCAvipld
VsBqVhEb++sf5BW8eBPtwrWQHNQ5Yf5IL3+Jyr7SaE6/mZuTQeBMAH4Rp7sSI4XNzFMg0ZQBBlnn
Gyl9vCAEtOVEosbL9OSQy5ZjJ7KNHqpkndatvn/VnM6BLcQ3Nbo77h/vqtYOBnuIUnFjHzpSPlRO
RO/wd7jQtA2XvErOKZYVobunIQcC20inKneOlmO9KdxzsF5lMCLuBQsCTv8SktOwqXq9m9RULs/h
cDgCPw0u22pgqRadkCByK7NPOhv5H+++ky4ThgIDZqIf9hUKROAQkJ9HCQClJjTmznw7zfZXEYpk
tCu07m3DTu0ytHfrM3f+XHRhuJzVzr0248DygWzhAQ6jZhKXw8fpeSKDzAhP20vvWQ9ssWt7iB4n
WMxonTXIzIpvnK5jO5vdrpUbiwIX61Ifwk7bxezaTxp/FwNmHMdG0m2mbRSs9uba+iOQfYl45s7f
/UmGuix+gpsdcAmY40PYS7JTLTwnZJm2UfVZFEQsqAuDLO/ON/jetg+DdXDKukvoOOBrErwcf2fY
6ROSfU8p5lwtA2Zow9FmZ2UGCP4k9PqWg6OhEd2DYK4T+lXEt6hhCEQ5EKtPQWSZbFcBqg3kaCZG
wIuMOoKoXRqrlhle4eUACPxTgyWNvhCC8KOyOhlE1EOp2G7e0FJNspaYepQ5egZvDzYo8vGVdxgb
wzrQBcYM3qo3f4zOG2NYMqRQllvoieYdDmsPGp3KyBurfnEA6ech471NxpOg+dJHBJO5kIe6srwi
o2XfPlkfEB3/DQLWbNCbUI1RKiMMN1TxWGw4FXJY3BBBtCBk5lO345Or8WbK78BjXsdpa2gZ2jv8
5PtApIO+6n5dHji6ODQ/PEe41iSHSy70QCEB0Tka7ZB+V5rZkgWxlrxdcxi4zKy9ynEQpN6AmW82
hKqJOXhHMT0Zy3Nc5l8pQxX50OW1Ccwn1a9euIr6DcYyveDdD8WxngBENk58uCEla15jyYfp/f6j
FFLG1OAyy2U7tQz4qupdd3CLg44A2lSOG2qZ41xZcDU//aE2lzcJ0BPz98J1F8/ypj1RQDeHV5CG
TEsheHQghOTjdRgnOD0cS0OM4MArW8082k+9jIrpJIHjYh7n8/+kBJNLgX7IkpMME7saYCzDkWtP
/r5aKBaFF4YG5OFmPNd2oa/sclXrbB/2B2i6UtfvdhUE3HGmURQICAQMA+DfpsinKGSsn1s22YQ4
L1dl/m3xb/lxb6xP29Dr+RRwGFBGtXp6sbhvSVO/qCNYD3y9oq0rvwLZVOjHaTUlag3xMHXD4TL5
eHOPMJ18EFql0GFWVk+egClVhLkPC8nohbv+/9f8lFjDtu7JiTIeY07fgu9Wn+xuPwBuTWk5pcax
2BwxG/22UrMXneTMeoks2ezbyhzd0bILRY+DqnUhASAreaB7BhnDPiwGKkIdq644R7PqHVme28HE
Efyu7VOFEswAI58AdsRZjPs0Cu+hLakmXzSSd+f/GnVup6pbdVqFB6My3L724KC70lHTCP5SQ3EK
wo1r/UVQsRpHOse6iomOa4W+Zdna/wo3K4QPWqumIM9E8MUCNFq+boGmcicjtvmjEQxKJ2G2Sekt
sBKXxICnZrTT4g8SXFrPymK/IYsd+UrrUA27KwapgdDZNsV3XlcpGM1OtJoXWFoy1LNzStP/B+yA
mR7xjZD32dJ9UOPUMcQRk6rN1p99fuB6z4Ww3UpEmBY/C6B7huth2O5h2YqPR5KggZKyHwXh9Uh1
ZI3yJYW/L6E30asfA0jBn3wykjGqvYhgxaL6TKuOeXtn06h7pE95MKNihqC5//f99kxk8P9OmM2F
TMYYUOwbW1w09ZJLnJva2hgI75SwMEjxrRT89GJxFTKt8pdNCnJCjiObAy+TE6ne1Glm2RZUTrKv
AH+Y0Zm/+SY7hKq0dX5B0vaPa7LWUn/1h9oCEWWES0lvoJqvM4LUX2FA2RtkVYjA1grNsK6smdvO
BmM3he3nKqYuDtyydU1xZ693G3liDUWXpKuUNsj2CTaLZ3LmaTeE3p9vvd6rw8nxoHW7S2INn5jf
J77Q3WeknclP8jLTK5Lhv25YD4bJmviF8pEQNYrGEzdb57lDz/A2IfCmXh8brqnCIe2TLtmKRwZL
Xb6WMstVsb11dYSz0ldNU5/6XAJSPU/pr0Ofzj1glbnNMvdsq++WILDBsTDdnz3DUHZnReNaTliD
6UxUenLimIbjFDae7cXIZwETnzWb36PFos00mO11Yf+1e9kc5Jbu1ZmAC0RsY+5avOEnyxTZ2bj/
i8a/Im8MTLA6LhSsoNXK5P0oEAIkDM1MhqoUfTv5jVGT0JYuXfdWAoRbdpSENx2bF1mUAcR1lEZh
Uh6Yl3wxSj7bPzVa1c1Ng7r9Nclc6Dkrr+hypE6JB+0pU89xChm7oFsl8K6kB5yxwikRFhAs/HSF
h/nJCD/bkOCMQtgj9yu6O7PGD9S6BbSNUBWEcyM/uHu5M1u7Rzy3Nboe+agSCfVBooJjnbQtDygW
MF8FYe1bZ+r8PzBtbfACGg8zuLayr4lJp5B9wv0p1+61HT/IDlx9NeYbF3h7dj+0/fpo0LeY8x4C
e6a44vEfqMZjqpxlGnB9VJ8vhG1GxOxncBvlykeedS93BxQQ3yYDxwU1bgyCUzekU639tAp74SnV
+FxksBQhpdJ7g8LO37Y9i2JYfc1srdERWUpYOQbFszBydKwEtHmce9xDSnL/nzS1M1dE/E3OkNVm
c6Qy7B7BvbwLHJi/1HnvgmAceo+x9WtuvsPsXzl9GE9YpGGRxtQ4xKHH+vDFgtj9G3yL6dhu89xe
lt7OP8oBrgjnSK61kNagprsgWuw0PWqLQU7JBDDAbq+bhy2IFrm3b4P9LBi/QiIJuJVYa3L9aCw+
Hh3VLmxOTwpwqt/kmmYqlnGqpnf27j8B+0GqT8wIp8s6qMrPLF5W4nbBrmhZFIiVfrjDgGcu51++
tIcWg0QhUX+vbASsoJmAtpsnT6yAtui37FxVBZCReJKjMr5kXHa9w+OaEF6xRyD0zgUQBY4FjNPV
0kcDdEdXA3R5P/SnrZfNDhCg4EylQ78Xi6RAWEPnyZPlpLEYgacxO86yWmD3+8jI2FxePDMSJfPD
qc436UlrltAGM1tm5nQv+ESxd2y7H1peIwVfkLjyFAsQ1kFTc4nwTVW4/VGJDt/fKnsjeKu6c4QZ
UcMkcUiKeeKLvoNBhShY7bT4U6Y+wnyY/hoxG/fSRNmrRcJG6rmJh7xWRmwxx3QxGcHQleV/tPq7
CoW7Ip+gT9K8cdvJXG6rudplnmSWSJxm+dv0o5i65qEXbmF2hjXQ0NU5ent1oQwDjZYRn7wqkbeA
tRb3V7WH1uNgfwotRlFLUU1+YlCgE2V++mOZdzTZJR4cacDtgekx6Cx+XsplJXAiFghDEoWqI/zW
RWEWlW6qbZ7uEndFICOe4yK0g5Nq9hyVeo388mXyQkEwu1K0/l4waRHlIACZYDqz9GfpFxG/eBr/
VyDLTepw8onNHKYF1QyKqcHF1fD/pjNgfT10+bR1gKUMi0+YzI24kjJcJpPs5jpuAiHM5pG0wzA5
/NNailPCBlTQ9GbKwwOrKMF0rEnbkhfY48z2xkS5gR9Dbe5mDAtxgEyXaobgbhJsYSWCLZ5nfSxL
ZtE12paNEZ4q0O6febrWqWfo+zYqbRV2qYZzZxE1PfHM5Uo6eLut778oTO98OYpai7MpT1SswDdl
Ba6cR7kCtzYdbleMPirYZ1iVi1+0ck/DqPkY84lYfvcQ139b3o8FVYHANv3+6kMx5A0t0YqJyiyC
5hXOi3MiXmQDz/hG0LHv5oOBhc2IXNOaJ4maK7oHViutPuOppEWIHxWMpHuZBoebNifmD/RMXyYP
eYr/0fb9mSwaPSSVjc9kysuLxtzRVxtZ0lXrgN500UsH5CPGcISQRiNBtmkxTQHLnrdlgXfdmnnt
tuamMnN+Y1mNqFfWXCPVlt1FCousoIhZT2uW8VFs74qfywlst+R5rLAKidoDxOOaWXk+eWwrJy4e
PTT/X6zyYqOhB2/kRdbsZwSx3orjB7s7sNh8+FIlkneFhtfOYnDibRIntBKd/TqAD88kppxPCF1h
SoA8mE5M4suaUgjaz9KU36cTYCY0sx7iT/2dbtsBUMDT4WXHi1u/iuj3lGPjZCxNy3c0eDWbGZeL
j/Ry8LG7cABg0+pFLfRO0DswaPIq2di7DIRwLtEnQpABDr1jgLDHiowIkocLLN+r7fWJe7Lyq+fu
kJOWO2qXbGSIKLKyRMH/NdmDpJbb+JqZJ00ITV8kfed2NrMYZVpLa/+FZtzFyNm1Gx/y9d1cqOD5
Qu5JjhngJsE0gCvEG75KveM1VhV+0kjq8wpHigAAzJhJt8vbFHStDnLu2HygydZcuSRZM6rfN+Lo
8n3WypeZsVSXApxnPB0Y9WdUfsPP+8A02S98ieLQKhfJ3bXdFxfA50uwqjyTJz0sjMAy3YhpS85V
0wV1TpsnhfPfK+wtkw96uqxul0otYocT1oa86Pdh/idwb6O45IUCXs+8cW4+utS0ZsdM/SXmEf2P
tx5HL3XrEuxFVlREF+S4sENy5pqAm3uHX3uRJHmPQUhQv6nUdqyJjbrnz2b03cKQribrXcLNxNxu
PgXcXwfDScXBPZe7l2xgncOQAyOc5gyevnH2KUtHdjgRi2qGqHBdrZIfGUzD2+YTYQnCd0pT7ZdD
QROwIQ9xSWa0yiePYVsBRvSf3VfNz3h6EIwinGrKhRSdFiTa+hf1+peetX8HVq63tL7n2eElVe/M
rT2epzlZw4PqXDmxOZwWgwxUGwk3jqC8aIYPHRwkdH6sXGlnNO7wOmGEvGFLGX3H314JNUINYGET
QbLmAjG1lgIHMJC23kDK9l0AZ8Tux2hkng1nkn6F8CUcaX4pULrPsANQASG7VPI2gv3ZEUu6PcTf
4UdP8fm6E7Yl/ApfUziwnwUAi2x+n7vx3V63lQdo0W8sIDT9KjpROunmIfZvqGMC9ZVBIeMSYtvL
DukwCVsIHVOTRBGb6mu1el0yLy6vahMMJK5bs0OdvXmPnJ6EhBxLO8kg/0PFvCWryOHs15s2LbWT
JE7q0eYtJvu5beyAPR5m4cwABw5b8loUHmouqvesKEEZeYhEVCo6qQYnIOgsjrNVvopFEmZ+3f+z
wt0BGjFKSRuSFZAXvM2nNVbu31PjtGUmzK84VbjyQ4MMfSixD6LlWX43j+eRSHhHdbhb6/Fiq4xd
ft1tQnjY7bOQbUFtWtNP5Gsm5IpkUGS1cSwR09YLiKmU73tw4Gd/s6KteD8RUvoaWTSUNUYNxKzD
Ecpch4JaPpmNroccltvtAdss+v/ans6zSpgJFLSy2Sebwi4b3f+j1KwNJwAS5KSxOgbDmLH39Rp2
WWOxfmOMasgHnmkcofZIxRIfSWLYa6i3RD3gqlNxLmZm+rbjB0OY3JxvcfzISMobTJrLoTfE//lU
78T55wV6Y98ILZeaiPSTHJeA9E2eIQq8H3EPO2obDd1sf9VYnusBQMg7uRQNEOJd0/e+m/tzsaCX
uWFoMONKZ8C43ShTcig3S346hCTWXRrR8KE/NKSlPj2OEouzrXpTl8U/g56/gQOuAn9EJIcu1XHJ
9L5SRGJJQdSBcaGJEQUFq+btn0SFKRU5EEYJCYY65AqzxvsF2NAvbYORf5GT7MG28v4DF1Htukpu
8t+QnCD+Av0jr7RLcZbjdj5iOzj/LCxFGOkBOgZvkD501no5TeaGfniag39cpeitWDFyOgRXHonM
OgwVmA17OrYRzDvYpHhBnZ0RO6cfWM1iZzFcC4Ui31rRYgUHQsMBKO5Lx+ccDqtRpLhYOmMzfw1A
5dfzHYmWR9/UE0s1wTzNn7oSOZ47GmCL8tYgIYK59KSz3Mowb5D+8cILRtqITR4CZOzIRmHBTMKL
NEdV61Y32M65YVLQ5wP95sDtzviIDM9xwXN9IcN2uvk1jMvcrx3/KJjfUDF5KUpGtlMNDvfDAbjh
pik4e6fifYcQCqflrQmSBRlzXeNya7N1PP4AoIQ2gLfeY+48Lyc8UzRu9ZK9w8qzpITekDqrQZiN
tD4Mfzp/Y7ufgc9WKy3+Acof5GYpQmb6Ws4UcmRjo5Oqd7Pm6rw+Ah4Uhqa9cSD+zxOo5Ih8Efov
79TmnNRwUCPwsx6Ny7zbvC7JdwXFqKncBipA18WmWrTVT+akgEkzt4si12gqVGP++5e/UEcHhZWX
/DriBKlsLmiX2oAr0NFnrZrdCtN4vWJho0Q2KXUMuHlR3qfKr3bks3MT/KimLf9KKW/aRo/Wj/w6
YaZOCEtcBnXDYbIUKUs5dOB3akRSie0HC9oDXidejbt1pwUuFqhxyCs/JipAFfK3F98QsqCKIcm/
jR2UFXGxzv4Fcn4rL5/cqv/ZO8VoS2AZcaFGnazCpGKgtkMTBPSbpr3sppBil4kqPcpAiRzAgYgM
Xnp0SjGYhHqvryktiOON0j+gO0xkPLG0BURWV63q31vw0SqhCG0mI+bZeaBrSYCzf2njiGbo4gtF
GgoY2TVwff6l0y4/TzYBsgPsMbogSgScEBqRB9WYawSc1l0fnvPbIapCi1fQOu5L4NVRkizbQ2ea
VZKYBFBj4867HUxi8DDhDCO0iW3vQvo4lpuoqObezMESbuf8dphcKGPdBr1KetvEekmT8PeMo0yo
Kklf6ccW+WAG3oLS8wZ/llJCnhj4878kaPw/Oe5IrcpweqONgPOZ9lFuLcY/GY6IFzzs1Uq4tx/p
VDGwwUC+5bJhzGV4WebtWfFhu1TvhpkkbVxgP3EArc9al0KimjcxLKErHbQIhph9uFD1xva3oAt0
m37CJujAqfqFyQqt72O7ClrMI0gmMD032WLjBAaDIIOqUlr54bkS84el1uPQ1gELQD7jdwMNAsYh
zo5atyYcLZySYyfrLK8aINnkWYEvC1RpZKei8C5y7mXzIeuewacMIzG6LRIllbDVzIXI7pmWcH60
wrPtTzfzxMkj115/utgMSWUsxjRgFLRaxhn/1ifmCqhvXoVT1TfLvVfgsy/+666a20LPzgMNqx6N
PKw46+5NNgTd81XhiR1HMolkRR0KlggSA8IZ5BJQwOMMzJgiuvROnkgqcnurSQkt5PwEHhTO8e9U
oUvTtiHTGJwdpNuTHTikwUmXzAv6q6ZROqBmdtauwwPBouqfpN9Qth45CPM3ghCZC+a2Que/8i7T
F9GJB57OgL3Iu+Sg8EXOkzx5Gc13xcbuDGC+GpPQlHoKxbPTP9f7oPvXbZ4L8uPwaZM+j3WnLJzB
f1XXerx5Tgq5jFgZCIm/BxrXDrH1GRNC6ZrNAYW00ESwl5cO3orr+CPiHI4mhBWxRE8vTGOt9FgT
T6keHxgSRn0n/oaiuaza+igMzcmUa/u49tDNwdUyuiwObvIaZii25x4kjOG91fOKoDztCQSvJoP4
C2CiqM8HSDsORycr2Jr6c4HA1ORu8vGdWeBZubspJsWJFaGU8vYposAiQdmoeGpshBsGAWxvXtEG
XUq5amLA42R/EE6V1XkqYLMXt1DNZQXObwY5w7aYmi3EWtl/syg9ZQ0/gRrFCREqWvRdA/SDsggw
pxJ//nXvGc8XVnLWFCtwJnXx4gQ85jOvJjgK3LRiKAhNFbOp5skHNGWlSCaHZgS0WnYV9bSp6Fbb
0XTCoNuha/e0QbJ1peWyjrxtv6DwO6uEU+f9sB+NFglUeBzBTWb5U26jHp7Z+hEshYB2lzd5H5pI
f0oYROLnN4bh6OuJuGqnmiwACoATNux0vCjv2pxeaeWsv7k7ypA0dCnlNB0yukyK8AqMxoPEsGwP
6x7wkWEV1ePbhAmJ4yeSPhpF+C3cFhbvMm/g6VCU4jZBjXgQqZB0RPUTnt3n4dKKTVNRxzVhh0kH
EfnF536AYtfBYmAfVFN1BmB1fjrBFAx+lm/HmQB1spbL0rqF8VaCxI6mrc7aNk936KlcnU2SI7tB
XyNa71RQE9TDeYJZNFsNkBdihPol6iFNRUgxTITzX6OICrZs47qtqzDBkq6KeE14uKvR5sgyg8cI
FrTNMc5MofnRNg/1wtETtf+s5+WVLlL6DP2rqHM2vkgfez3LIiRmi3ujayrEqBdK4YL8IaV9o4IG
ICAbzmSTyTCH6DlV3cYYll2k+cY1SbY+Iv/2RPJXCC7SgT6CjSbUZu8QHGNJ1QsA0k9gyowClwjN
7BrAc1uUC2q7BQGhCKtGUCFXQuHLSEId9Uyu2QaZM/Mc+ElsVDzhVkTvFYCgtmYsNXruIu6TPcIk
o7ZJTn2/7YmbsSOkaxpRDM3EZCcBOVG2QEUYXU+LFdmbn2BpxEeEnJs9zcYK8jliFXRGVNqS5C5A
3iYozgpOypd5HMhH+a9GrIiH2uacHCLYS39AguV+8F/Kqku50/c3auVztCILBL+T6rHhHEGgjKKs
YAqiqztFmqYSxIQ5KItQJBBn4/xV7pW4Cj5IvO9UE93zKP5s6eu4jEiPMr2X04LaP+qF48yV8e73
OsKL709Hax7VOKY9lWOoZQMy29WTLNZc6WpNxU8PKk7jFlckQkx9yJSGxXu37YaHWdsx2JBpV+2J
LRMbR0m/EZDZJ/k9MkaPK719ZwVs8IWH69NW2xBqVJBwE7oko8/Az6tWydHFdCKjc6JBC0L5r8zV
ECvoRytGIaT0Oq0op/OII+jV/gR1neS9B7pK5QeDgzou1aD0HsObka973DZpp47QaEIBZ4cyqO/d
ONIp7OO5d+TW2sdwVPmu57hw7w01tRDxXQGuHBJvAKK2O6Nf9PDTEbhm5Uk2i2NQCwJCr+JarCAp
KwOVzwNFzkEXzX8VzBTcUhPoSWdR7+dSd5i9Y3f5/I60xhaO2AfIzaL+6VAdWdPiGOFQmgTsHLmt
Q76DMEttizxY+Fge6qzpXxSBMVZ72W6q3Ofe4Y/WawGE3JzBMGGS3asyei6IWOoSMrhzgTbzWPiM
dzrATpv1pdLdX9QIx/a1RIwORuzfRL5Nw1CtsAJaPK/FtPzjlb0gyyQw0n358ohtD+louEjZ1FEg
zLrJp1+6YwERKVr2E1FTGxBDKuAklCVHENc7l0cr1U5Tzs5a+XtvEdP0T1O+KcUGvvaoFJ5VcZja
xrMU1PWXKzlkzfsbWGe6LsQgTIsPwu4ZOrVCqZ4UhQw2uDsDf8k9TluhNWJXgr2uT9uNeQx4vmgm
MijgX62CtWdI2I6Rq4m0iVndCvpViReWX1H0kidaoKcG7/AVhwK786WeDRk23HqkGKMVKjZDmHJN
ulgyPf/4bPMk2PqxP4a2rANPMEgdYEgSMe931CgVUejBe73dsJG+mZiblDi6kKmE1KpQBUrHInUs
vvgiXrtMEP9sVHRL2reoboexKkinAwvK73/hoM7BMdbRvD9wybUOygBFsMyyQyZBrD600X6sOawm
QlP+wsxfKNi6yQuaDYxh6NpaHJHPPygfGuMhjE8FhTG2jnydHVo6MpWw8EYqGSaA4IOl+T1vhLgN
UCLOndss+wlgagbNcKuf0siFbRu415E4xO+XFYTVlfgqcJFVy989ErhD8KB8db/aVdKV2Hb60oll
ZiZjqZWmPaXOpMgaHqazryLYQq7BbNCeKOeIj0FlLswWuoUnjQ8wbI47T1qgot6VvpGZ57HyzF3H
/+Bx8QKdhxNinDf8uOkDXgG40yLU6nUpQgpRmjNhS1F0yZ5kwYR68CtCELFU+KW6Esx2+lYPjHr4
CH6B9Qgz5REMbFkvyalm9uA9b2Ixc5Xb9oMjUL9H3ATqVUBFuzoQWW/Q+mN8cm/d+GZtxWk8iLOT
Gs5SUofFdjpRWwvgRUBFOuGUAy/bdcEXd9H5bJDnFtGc8x46D4tbecRU95aC9aG3zU2vHHbuZD7k
KXxgl4DZeSn7Qu4FrXVzrL0IQEhFvB10qEyWgOUayx2m+GoHjKlAiaeCSL/fb0ppSTzMOvCK675F
T6/Gg6pZzk9puUyoa7sXGFiI4ILWRIlqp70DGW63heDaNnyfnkOiJepgH1XS6i5VMDV9itXnMurO
coaUyrzFnj/mohOF2AAY5Kb6xrL1kyRs8iJ20YRZmFylRpLdYC2XXtyQaCk19YhUEn503ACmaDVG
c0H4HdLA0C0SR8dhcsi2RKugynWVqXi+SU6LJjNGby3FyFtwKtukI3LYYUT2LC3JOJVBIdHXiow/
KRtrtCH6VWA9DOUHKohPgG41GQoOIMbX3EWPbOVsO9BLJmSd58jINtj/kuIsOcwZ6DTvSTf02fQh
aFVrELdNzP/npwyz2CUe6SVVehGb8Fb1vXmasVDB9+qMN5FewMw/AQ2bOjityPKQncos5mDcZ8LT
QH8Wq7N5RxYp2V/3tnJqJVsvuxrT3s1fH//bLDLm1BbSiVyC1hfdwW18SVA1FPkemh57Hie6bKiA
Q9aSQfpa42DhbftZllVfEy5xkB8wfkX7MaFoFCn8uJQEew/xv9PfQBk2OjITIV4rYyuj+VeYJGdL
p7g5qTJnyE9pMXUBdX8RyA+4v5orsg5IXVczX3u5sbE4V4Op9ePsOsmULScrH3gfBAMsctr7KA7f
mxAy6XCN6J5mWgu6M470xIkavpcy6V+8RbR9y7VgFw5J4NU10X1zoIvhIadQIL+AA4ZWoPyQBiaI
PwsPokPaEzAPKMdYN4sPvNVqHZFlAU3ian7s7+qsEdMadfg13JcB8rvm7kEjWA3kW93p+YSdAhKI
rvtd/J5kmjOnQWNsy4HZvVeyI/Y/RAFkv1e09Nn/rQ97d5378s0+GhDzKaCFVHVRWSt4IZIvJrxo
QE0QxyjDLRaNahonMduJAqSDG/ibGVmWs+GKxPLY5xvLrd8TR57BK7hPDzKia03eDASLB2IUdE5j
C5eVAuISG6xPnURAOaWWJ6YIYXHIIX09AIRZWGX7EAcR25pkznBmrWvD53mIsBfCGFsTrXjenlYL
r3QZeXDIDOCmw7q9aDecTHShZsCj0mfOt4wxKfzl7sBSRrOVae5OYDSWDnmMYJhDKXDpRL3vzmSe
4U9KFOfLwPjqh0ZOPqcr4ICEBSfWoweWikAPt/jID71Eh+LO4h3DOrpU12uF+YK0M4k1jqrsiNnC
WGonMIIvpqYknfuVAvcZDvbswRJYXnSqZFtGy4w1l9McWZWTrGT4atUdgaSksKDeW/3U3lft65UE
o1Xvz/Rj76vaV1vb4WmoIm6ZT631VMoUtN2urNNY9lw0tvXUpyldE4r5mzJRroKNXuYIHHiE7c2r
zdOPLYDkrf918hdGWkU8H8ldkV8vPD76/m53RCXBYDSBtABj15OSm9drX4Vwt2ilml6JRXloyy5f
cMH6kSy4txzukwUG5ReP+OjVAi6JMmrn0yQowXy/CwHVmUrShi/QMfhBXhH6zidL4+kdWiGlI6Nk
AQsvG2E/LKrg9YIJZ6RmoHo94/yTO6F7EXk61ZjlrqITmmQ63gIemFkI7YgWD1kKUNpZGQWQLfBG
oN/VlDjRAoaoZRAy+glRj1bh5kcsHWEEoxFlIE7mDq/ehEUqtYoLsGPLB32d4Vq032PJPLnBNFrU
YvEtdz2oGISYP/OezvKy1pApgd8DLUnFA9/PhtePFeADdh0fMyKRgxcSb6wuelRkHvtIQNVsUn1r
Onii4HoicjeY3zZNLgx1cP2mir2OSOiUz7Iv/EFpfBcFoCK/TFTkV9ke4KFJTIjuD5ylQNkL/3CX
3B6hB8dPZr40WIuAAkkcyotrxUSB3tg8g52Afewxk1Xu0awffINK8VHgzkrgKxyp+d2urPy3Km01
OPPR6phVW5otPS/U0KkYSJIq8w04JK1mcU4kzQ8TW1Ubk57ruWJp6e/OyKCE1F28QDdsSUQFHLht
l62+jpdy8P3BY1pE5Pn8/wy9IaMqsHrxMOazM5bZtaJ3wD85hnAEYwYf3AEWupgtxkMq7WKjuCUJ
Er9Urkqo5vQVeFzcq07K3zBMNSpbzXpQvkzQe9snp2CVFXXGfTdKr+woyFZ/3hZUPqrsnndSDSy4
yDSwwUV1uMVcaZc7rUqk6QaM8iCsTHOc6M7S1pLv4soJxeUp4ecxa/2rlXeWIiCHQRtcSiMhi8yL
611mRxdpVwIgwrikzz2JUMT/oH0G3q5k8Kt2ES11Lcur6x7OImYq0mFpzxjh23dVnHC1Cpp+xQNJ
yZEmexbjUrvSNgu9MOAfHidw1H3ztfgGyrRfzO3x1GQX9Pk/rSjraU7motgEssns6YZQRBReE5aG
GQD1XOGsiSq6VLkwyxuYWvrV94UqlVCUKqDQHNKwjBQH36UPKKNgSOiebIpGyGx/e1EWZpfyXUkr
+k9gEjfUcrEJNwSlfx/zgtd/xkwlYCBD3ZOkRzoVFudcBIzLol/8QSnQ11KfXoC6cZPty1DR8rhG
gX6J+A+zdHM+jHnR3LAch5a4VTbhOAndNozsFD5p3bdhn/OUWyXvalhYBD6/OLXsd/DV/UDom9X6
DUo//ntaat/UtT07N5j+0vkxgibBL3CdB2EQn5GNUXZb5peG3PJ1jdGIzGMCv+iu4mZXWuLMPqj5
z3ruI92JER/M+IPA4XAMYdLRoCOi1LPQAI/9phAloLC1Kvlfa3bnQ1qRPV8/lh6BMMN7eCRHu6M3
/YCgP5x0aYFkAb5s7SnFlQxvRMleMiGMIYXO64Nc1/dRnxwKyvt+xcWgX2yYsK+p5gpTdwkS27WH
LJQrzfKzGFWxeFlTgdBOktbslLNFbaLV3kd0ocNG8sYNSp/OZMbdPIEcABcQVtDQ5+bZ/W/5m2c3
vdnaLMVI2DDgojy/sICAuyu3kmumAJpB/PaxlBWxWh2cPfivErLLSSJr5Z/W9zsabNJvzLSB/DzL
jUH+v5yN8W5Re7sQKlWmQwdqTgHO8AeBzhrTZv8LyYnEAw1aG0hAjLwqbLygHvtqmRBBwSLdsJan
QKXCoaU1kKVfXKLvHi1koLPc4DMrTr5CiH9QZHtQxL0aZhxQnwDObFiD19YLX9zzaO09A+S0QBCF
UH70rtb7QrFuCP+T9hmsldJkFlwf9gIQT8qeXwLPG3ep8Oz64cACjDsv8BJtNqv1bUKZEFSiFHaV
V3CRGpTIg8t7TsbqAKosc5SAKKQFpikBZ+gD1GoGUM33i9sl2VeWqLKZP62g5shCpacp7ueCH7wi
clZRvys7hBxCzwznS3GuYzFIt53QrE2K67I8sM/4L8ZVLrUoDM+saS+LumXWk+ImmS57RFQKXLM1
AkROVgL18KqzUTN/VDQfXX+9qHlfL+P9UY/VJr3XiStBr3HnUPd4sCo6h+Sal1RkZZZsTLMSNbtT
1+pnfsX9eL47FJiXxoX9nwWWL2AXfNwUM61F3n92X23c+mYtUgUwwBroYwkNGCsfCHcGgDtPOizh
a+eMKFHb+LXiaKApaouu55ZNAvJ0XyV2AA06lAMsUzlRH2qSZrQhCuwxlWKnaBV/xiNi/pqMJ90t
tBwnI8bKt6Vri+Wz3O5R7ZXs8EZEjbTD2msCmAjAAGdA7NhAeDVZcGTukdytjtsXxm01q3/QEH4A
ChQ4Ur5jhZbkZqt2F9iAoUiVLWyivq8TubWka9LExlv0fw3Wb75CTYZCWG8fUoKQYARX7tF220ey
ukOSS7jCLYD25b8ESNxFl7ohpW6ALeUQ/qIBUQTdEbx+e1N2/FCmLS7VFl4xJ6Vc1WYgQIXylxWc
xPqqLVY3nLkoJMcJ671VCD+KYocb89IwMoSYQhVAkfHRXqBGc4nvrriKwOyr2IqriV+Vp9KuPdXR
roPzpAoY4E/kW4yT5ziLGTskrH5hOyPTNMUSh45tN0KuzdMec0KHyTQ9fHJuZ+jdkfu8G+TSIaXq
Nffq5qsYPzxppAmb29p0hlCupnewqbVS8OHdKAfsh1kF1ekdZ6bE2LMEbXGxEZOdY+DqikYwoKUO
alA6ojPr9SOtc6Ir9KgMiQnVk9uRaiAe1V4SSOoUsJvbRoG44LXIsczvV0dyWalYkRzroty62cPV
dDo8VZf4sywXp2EwJge59wKTrmcuGoUgKciNg/Y+Dhx7pinHsBIhm5ol5iVz0YlycSyR2kufsTeF
dDw4QfWXaeLAu7Bo7dVRnnc8WsSVBTqJZT6DuKyhT2of6cjqSuKQ26qRcw/cUuXf5bwTHnmgghLk
JQtAoQRPPADA9vM0QwTxyZSX68FwXxXG0g3xXWaS1COU3OqqfCxKedXbjDFeSAJfLL4kXhc34BmL
n5jsYHWDERzCkHJGvEcoLeukghWhDHuy22s0bDne33XCAf+eVMC/C41uS0oSYsvfHA9YLj8M3f5j
K9rLVrA+4aHrjWiwZ/M8q4S5Icn1bu/ZAGSL89JfPXZJF385U2ZdyeI72CYyvNI0LUMI3M7nUX+C
kj5ZvTnISkBZTHLAGZMPXq3mTUG467UdMgTKae6OYWJyaf7UmAJjzyOBji+crSSXDJ85d58UA6T0
MVSCIaKUKMScmZl4phWFglsnS0KP3JH4eiUsDxtSlHOtZsrh59tIyu2gj6kLF2ITNzMsVschEJPC
TrPvS+JJMde2H08fzeyNHJYab71/Dw6fIhHArPEhlgip87L1RGOSUZuqCltpgJyviAdSzjXb6Wsw
06OJDf2ucucnIS+/aGbv3QbBaFPaVeXOdqqbF52LuAbG5IenHj5ZjMPKIYPVJyKM3Ca2UnAwW1Zi
ccIUHg/xJV0vz/YeZanXNMDtNZX+82MkDS8DmXxXplZPBDA08AjxR3BvlQcdEnfWa8EW4GzTy1LU
Nex23fbZp215xpcDxIK2O58/fSjB83lNiCw/FSuIgRfj5n59uzi/svYsugjpfWGlPQpkg46UZYnQ
0WdqS5vvQ5BjwtTvbGBo+TpgEgjp56f7v3vo4clF5dUsXd89SX3fq/ct89MEangemN/U4eXCsLU6
exkDrqQ5hgjYy8ZmhprubA/FYjnQknOWee98xUVqnozi3NI14fOem1yNcGewJQmncH5Q4C1KmrfA
260t2z19L7zFl7PE8jfshRF3pITBYyeZLoe/xhq4UietG1+w/u8LoZ+Cy5937cpz20ZiWunY7hd7
hvWoFGCT5S0FmWywB8iue6jE7dpotIx+uOGJj5Xg/UNgZJQxBy/nSf1k0DKV5aOnIei4JvvY6Fdx
LjTegX4GmSq1nFMEQom5eNb2clViwZFaEo9GrbjiXKh0MyCfAIfLaDhpiCPIaZpXUQYwIo5vvDH+
9ahVZNOXvxEWmkE6Nm1aPLL4do7klYD4rhr3fdOZyoImP5NqStNh8eJFKODSw1jMJPVOEBZGH1Pm
H6UjRw2LKEbNDjHX1zlzOexKP+1ojGteEceEeCNfM64MXfyP4H1ZyNY3jhWR7joRTCXkWA7XvQmE
FCii4CcMKELbxhUhuqegrAbKQztA+lirhKhH2+9NwY2vKjmm9R76APdCoHpl44huylIyoJ0LZpSq
M9KKrdxiPQQ4fkllOiLopOEMUF3qz59FfreQ6Tb/iSqHSPqa2lLza1lpDt2ZafFo/E5zOEZEkLIt
IvuvysQAIVgm4PDIQZbO13Q4B14aFwJ2USbRAmxlkfB4rid1TEBI/GuFV5Cn7JB/6ZkiqVMvy0h2
yqXienBpWHtdwawpvJHxPuHSU2MkEbXa+FoSxkIUWROjoz9l9D41fV3J3AwE1Ar+OC7vS9vvc1/5
nEUjLg68tT/gUTHW1rb6UZFVwmNG+H3+FQUNd+v4fx52L3M3p6PRxN2XXiDrwRWiHlXHMwKL0HM/
XHc4i4Ztji8ywqNNKOFGHCcExB8f1P6rSwWcwC7KH08l55ItkL7MhswCsk4pmCn+UocTPvUdfdBu
Yv/SePB+4aWaKx10YlkCswoSmQsYu2fkcy+6wqDqkimaOkKc+tuKfca2LKylnuShuROIfh9CD5rg
/0AFIZUKFB4NKNjM3ueO5bS/GxAowrhD6OvIjdFJv19i/YFBkTIlegFeCSqRAYIYElkl67UvaNIq
IYv+Y2ChWxBlAkGqRwsRRgt0wS2MKLnA4wNG7bKvM1+ssDG78yKrW16dJjVbIyhLZMtBNI/O8ncv
Uyo6NfgRhj/Va0RH5inUa2uD4OWJZMo3IhlT2zgJ9avnxT/2NQ5gaQn7jqBDFTBB7c0glwGndIX+
v+baFxZbOoUtfg9vPcliUpqbCcyGkVnUqd+mW31Ku3DqsMy4y+D6saHxpaOqrlSls4FabKbV6Tpi
rS2x9v8PJvW43AGBZF5ivmpT1J7r4lwQmaTIjO8nSv+PTDntMJaoEAN7VDzr16TrpIDnHEQN2R3c
2AOULggx8no9ad9gBYIn9YwHUP55KyYR/3YMFgsEl1IAzHcyYXHXkEn6+w8WWDVbsaxZnZ14KciG
Ax66bAiAUvNqe/4/VvwJRA8VgYtmAfYzqLQvmmnqkEajvVR2bXZoO1FmHaiZ7vLyywBFDjFY0KHU
Qg9hLiP7+TuZ0OfT9YXATf+oUZII3kx4sMHN3f8gcnAczm6NpbULwLSfJvXigCTIWmBeGJ3NTOxI
l/Vs16EoJMgOg2iYGhiDV0BnI8HyefEFZ+WMmtOka5t4/QRD6VWKwB+VmlSovUEUghET0+M0NmW8
tFpxPWhK4/NwWeJeBoJR8AU6MU3etStaR/4ciBKlGcjVeBzzB4f+Me5WuhpIvnxOqQ7AuVz4PIHw
VV9Dm6QDXgJpWaPr/Rebf7K744+FiQ25P/+RbRc1qnhuVfzukSbRX7XTlRRZbzuK9RX5uuHUQfkI
eSDWKOfq5Ktj8P9Yq37xVr3q0g/ALmySPsyKtF/I56rOmG43WQuT1+5rm8KMZyVyLAHWsHneroKp
gqPA2KVAwJ06h6kzGjHBOOxQLYVoXPiH8EH0lv1h8Cq8ClAAyRHFUf9jdpUWGuYbPtMkk2SjOpo7
M9tXNMgpfuUPlITw2TFyOqHc5ZffVjL9v70Xish8+p8+PWT9NyUhqj/E4GkpCY//pQS5Gyo/FcgL
WMXUTCta8gaFuz+A569lhBRw6eo6npcgWicFKIgFXF5XQj4TRNywDe3yJNcUYnd2N79jCoodivG4
csoHVyEqXUgzH9fDdh/WiEjKibwwkrggjvz80JCwf9o6AN9nbo8sXzakrG9E3Mj5eRp6dl4ZqAed
HO1oSkh71xMBE+Proxw4HoKV9wUnfhxV5KWK814IYELmHG6pQdOY52eqF7Wk9NGgazh7qqN4cK8L
Irz3ZdDl0BohJ+spbyz3LwSrOB65ga52MJoKQ0rbezQl/ygn8ahXU2Ry7iwp5zHdLT8TE7DbEObs
YQiKNkXtL0ByNUwBewAN3cQ9wa1VYO4M8jE/3qEFQbhuHPhrLN/QnImtY+CZfUE4j84Ie2dk6GSk
yGU60+/Oh/tR4n3ONRPGxvK9lyY/KEQ3eNvqCB6V+bDcp4o8L1nvmhpgnLVEKVKVqCMucA0LHLPM
5G0SYQ4ZT2T7eSMs3fof5kGsJ6QsdYUTQaecG80TkUQZBirBlWSrN+05wgr8fN77mwUZJTPunTJ1
t7lLquF6l8kxdtbGyhsAzN1iRKsBgi4KIWtfJ8PzW7BkGN+uZsrIDNKlpoSVQVLvAuPUQSYp/ZGs
yDcw78gabuixdiNHN3oZYK6Mw40SxnBzPBIxUngjZEPK9gx2N3AnBWuqZYCHVM9P7M36YZc1QZOh
y2ykvvyEm/c23Q2Rue2BJ3qVzAKhWsiKeS+MiVMyRDEsRJl48RQo+2MMxFwT/19FXxiF12w0FyRv
agGVzIGMYQ55FPoyLDo4YPPuAfn5Dl48geF6hbg8IW804SSqc291uqT41rjneEKzyeTvH1gOHxpX
aTNnj9BM78BFmXBXiT0EcmzolQo2J1vXy7QB6q1FPUmEqDO0TIOarclTiok2lWu49qCvjd6b+MTk
hFxbncqvr8EIBy0s0zcd1pJbTTU8dAQ5SDMKBMnQClVd+D/AhcxLUg7GYe0bEA6eha5wQEtvcwD1
ZnJ8CaT6JVPumZ2i3pjeB/X706mVI22qL/0b8kP+fhdPabQVaRAAL5DcdFW+nQpC5HbZrF/Dyzw1
XIPAvA7RHGicHFawLStPv4rVpgWf6Silks5Oj6xPcJ52Welo/qtlPCEoulC+ULL2oIWArtqLWQ4A
h0/uKNDetoeR9eLANhE2m2nBPUDC/4k099jCPzyUTfdszYjqutgMAytfero59vaSiCRyC3SmMLU9
uIDmie+NXjXWUUK2Klq0S96JXq5SKZtnHfZ/UKfG/MuB+RCdJ3LcKbZbzonEJhDWxo6ttlUjCWc3
MogLkezx0Z9NGmhhpaZNljDyTJmHV/tLsUpXR5kD1sAIG1dLVZ1+pgibPHINNmapA68/KRJ+OFdi
29pcygVe55MdzlaKOBIqW4y9jNBC2ls8K8OXB42B5ZNlfWPJc+MAt9d9UybYF5txQ0blXZPD/+kv
SqUNnMSQZJkTXoOupw9eQF6Ku+rSb+2AdYaJiMex6F8j16pN1rWflCtuNZvJxtosqZx5LWX0LXxP
67aFHyUwPXE3Ofn64GBQO68xlpvUKwZ77ZsoXU6JSndRdOe69wHH+KFiBaZ7ZrWB/DWycY7sDhAC
o9+R6KFysAfbFwwskM1MKBk+upD9uPru2gISLfdquW7S4qPBmQu5g36hcq8NqYGfcgVJHJjTHrhR
9MuAPC+xWDptoKCZhGXq24e6/j8bOFSs99HNAepzYtCprOhcvT4kplxOkcmloHquK+6XU4RlfdK7
28za6oosQIr5mWD9BXb5b1urxOqa3X0kSOae+pQtn+BVDxo1lqcWKMgyqzbq4P+PW4MyfKNyTgVA
ztHVOVt/uK9CjkHZbJwTtl7KB5xoLIO60cPiMc5KHgXNX8ojctAYumm6T9CViMXOS4/hrQ3zrcM6
VuGQ96f8bnco2tltZvpb4bMnRG8RXGe+htBLx5F2sgeTil72PYL+rgCpdcooohWCXSpShmTDnimB
Uzj3nfC3YrLhi2IB3r/PBBpRV+WAySnm/G98VR+vHb1MzLUSKlSE+ffz2Z8YSc5ietb2itU1vcop
mY9RUHrgmzVl3+Gu8Q3sp4YrNEMC2XcsPhJ1U+Z3HJoJ2pD4rpFINetrVECxCCEoqVLc/1S0wMdt
8ufU4I1Mtd++hpFqCxPnxEKl2GOOmvMFNNLscOvaEb/ZXBloTMdgd3xEUoB4oWEdO69umTZE6Y4C
NDpeMNcDNnP4fF3lLhdU6YqeXIAgcie9ulxikRFdWreMrWaVR8DMMteNJaOKxDdRG9U34iYm6YT6
pdVYYmRyWz1TFoTiJxCZ3q2djxngFuh4zER2MOAG+Vm4HyPKRy8+BEdOoaT5jbpSWspdxFskACwF
lGOXioQvlFmHXyKUShNwtECAgzJTWtDwv1g2lWWCulZ2HnvBBDpx6jeLOYU1j3dp4nbHEB7y4BpJ
u1tpNqA801OcYM4p/FmoV2VVsBYBDqOcYqHdf+utIVKQzmsligpXEfHIS8Cb8xGfbx4oALGpUzas
emtOmkm815xYlFO3nzMbox+Cj8ngq0z4TGRILHZWcrMfrOgDd2bKXRFmDX6ZE3VKmnyuJlUa6Rmn
XPI7pKjVVTNoC7LXJLBuZWN3BpCoM6sCbHBsezJqjJQdagFJhdKc2YwpTMrYNHqrI6g30LghjPhx
1aG1/jOI1AjgJOnfKEz1D4ftTOpfSA2nM+gZ/HlfgvTurDJgZcrGZ8A8bQvFVMztLtkiPD0t9pef
kH8ZYt6EpDWoIjQSG9vBPlFuCc1igKsAZM6LXi1a28+jh8sRNGf2vqQfTSO4lB5fdKSPgQ/iFcxG
sJtG/LbjSqD2erOWpDPu0BoACSKY56TqdX54O4y8dDTyPOxbLWyEb/R0cRNFwEhTwMf6jq+iGkUg
Jo8FszTT8m6uwK4LjprM/UyYQiEQNbKJJE1f490ExEzv3Ry1snhbmgcXVwo4bEQJRoyVbo+C+rdY
rbefQOEp/nO7yJZFgx7yNlqJCZa/xIWg5AskKXW87XT7bJcedD/SXuDg4idHa6ekqZJJ4iweg4dx
UZYt2kB4X8Ik+JOrUB2gu5/PKgP1NTDyuGD/XF0SLqoKck7dl61fevQqVjZortg5j8WeVR003nTN
xZY9kHQ+0Wo+FaPBOrAKITLvw60sxR1G1ZDZglG4Irf06xsGNktljSw+FCu/YDXZ7icSoWERfNe8
U95rusUo/YZlgo/RbWFKM7L0WVN4kUkF99rf1inoa92V85zssgsutkIvBjphY22AA/yj3bE/Mb5r
xPL+YzsQIf1pa3xFsauFxsd2yS5CszwiZ+WZl8CQSFWX5+fFO4JCIVjVETAgj9WcJeYaHl+Ry3yj
ivJDoDRLf62UVpeXqa/WEymuEeJaBRHxoJyYZMoJLFAlxxXcEAl3p3HacEmTshabVQxqORB6CGct
gfAPmFBeEGmm4SNGHUU15+LoROHtDB5wucPtyirGqmcCA/XL0uC4Idy25NazUcjOw4n2Kk25l4E4
QGqSTBQ/MY0iz5UskpXQk9yZR59MkggEuKEM757FpyMfna+7Jo1KAz1wW6KwV2Z4+BusfVQVy+BZ
4F6hTUHlfvXYdc6Pf2xn/GTT/cVOwGZghLjD4Z4tdxasnlPn8pYppRjEVXGGGNKX4IAj1XZapc7u
rJ5baaBj8f4pvB3ke49ZdpEMQinjEDbU1Ww8vRVab9K2vxV6cxEQ8dwdqLksa0jaa/JGF5uI4Xtm
T9W5jofsDfe6YTYBTFeqqEGfx+9O31oUufCRnLvMJfs78Z/FV4TTMpaprN8+AWldfikn1KmFpy33
vijIRqXEh1EZjsuh8C2jhzVMJBZz9Sd8Lt63uzGSeopDnn1WB/IAQDuCVRSZhlkr2t0QpZUIR4v6
pxkRFw+or5m3Ljpf1jrKB90+JKPjm7lU35GwdPROCIyIwTJLJEEQE0++hr8WhvgCkaGTLWd4euVY
+RZZt23+hHnS8E2cPDnjtpyHij06J/wPRWf8E6H8d/n/AnMEpPb5fe3X+i608GiVhg9z23nGDr/6
V8IG/Vc5qMOvlyRWYA7FAUONl170/mjCTlmCLf3/8w5stG/PTFnm8NAoqlWPCJnfOKUri7U53XK1
n1JGTDeKzzPTtCru+Jk05cfHbFU1zE8UE/huElyv1VWKVrhtgdTAAaS/50R4opuo1tdINh7Bmntx
7NQCGYMTmkB72gqT7xs2sT0YVi0im9oEp+LD2sUlJkNHBJ6Oj2arkMiYGoAxWagx902uqH4GsZB8
gKcbto+DVUa82E0ss57rvsWQcPthNtjIGf66+0fVq3dE0bD+hnNnSantCbsvTDnEEmPWLTruyoPM
L/1Z7czFxV01DRjHgK2Ysk7ZHel4CR1zEeenOZwnW50vfLeSqhDrpfAmZZqvSfzFa4WwC7OpEXqE
l9nr+yxIp7hS2ZuCLGShdw4cfH0+Mg7dJTap9aDjEgy2R3EsyivxnSSwXYLlXP4pI5gcXhbj2vs1
clOPnYYSzWxvK2mFq59umUjNkKOdnWo71fu1b3KyXeAK5LLRlikC5gbbo6nNzmfAGQV+qGMytJJf
HWKbiwIJD11a9PtO5g0/kpPPKFFiOLan05BuMO17TOpiek5Jc6GyL8lfeRgheib2X7Pl9A5pMyBh
M8cB++ou4yazt531Mb5/vYce4lAw6VJnwmJDEVckRw9QhF9eAhx8lVbuFLLSLGy6mAP+/LgQDVQs
vf2fVOiZpMaGLcHSVLVrkj4014jYRYc78tMuWlA3TmRT9qOgEiqkizqXReK+IN6YS+e/Hx5LycB1
/y+mpkgVRwxf0Ob9ZMa1b76OeyrerHRajjNI2/bb9/N6naTmtojX2Y6Pvzra7LA5P+pdNYZfIxuv
RUTpxcI/2U2zL24TM8Pv5rZHMxlx9TSgO0Yh4ktBibWvc5TPum3NtcF1f9+iR2j3FzekX+PfhBFl
D8TYHc02HsKsMxgSuJnNKXMvvjEDcnYLXQfV3R0SfZKf7MLXqwMFR3xVTYmr9lRzENwBrJ6BeeRp
7+afpzJOd/5BXgWMbAxBwUNgL0rlbY9FasLo/Lx6MSNTotcUZh9mLpL494AFngO3HN2LtNv9aTFx
q8/h9yevaSvM57O5lBK9nkV0Bi0Q3Kh9sNrySz+NyWNLtAXS1vrImqMK3NibGXFFzYXT+tzIVmx8
vMzj3C7vGBl3wyNrRgNdXkJXDkXdxKJ6BvmDDXM2E3aCQxw37mlCOLSmosFoALZMn3MXD7ULee6c
tGCuMV/yZqgvcvQtiBlICPkETIm4FmJ1f9hpzoOn0dgvJajuAnXFmTg6AV4Ud7YMGiCfJtvD6nHw
O/MYNNB7i7raSyvcvzFhRaUgrdfFp8lnFE6h/lCCxg/KN8K3yg76HG54gny/Q9/chzTu/IRTIjz2
tdjlcQRvTkLLR2PUu+Zz7DwCCI0HVY0zh/EdRu4XTnX+hqSwJ3Sl7reK3dmsnhuiFcJ7WBsWLKyz
jIoocmHm2/nryAie64e27m4B7nAf8s2x5ehlXFRXcVA8BVlP7wGyl3ynLdnK95p9c0KsuyLwyQat
pM1nFH8tkwX2IM6JZ7yvy+6LMBcM1pTORuq5fTuf43fH6WQbM0rp6yv7wrValx+tWp6BR7iFEmrF
xNKpKb4y5KV67QTnKUFAy/WgBOWPZ2WPoHt+ce9nSOIe3z/1mpazkFJpyCH/iW3UtGqjKBARf5j7
u944nMVja9pj7dUIc2qT8/UaNZIOvxyIMRhKzvQiKVCgzXjjwgNeQfbUwXSXyYt2nFuNTBJEkUe8
8YvsOna/yXPRfGkixeJ2LMwuW4GXLEp6AFDHnA34y5fLdDrC7kiyLP7OC5Xz4HLG3/bbG0YVfOe1
DnK5XLl+lf3QYuWCII0qMVQY1G3/ws1h5e1tZWuMvCMrfqBnHguJ68giPz9eaHmPNr3n1uys4YLr
L1NVFPLDAMkpb/IG418cuU8R2KKeIa2HrPRzbo79stVoHOIPTzsC3ph6A+u8iX3Sy/61BqFMWryc
T5z2+orFgld4pwytdVkwtH5wuj2auLa6wNGG8c2tQFlbuxNzAjOFZAKa8hWeUcXNCZYLhmY7EFMj
bvhLT8Kr5zuoE1bM8gLmhAi5aiZTgmxTaOt2h46Z4p7Tb3C3W9icVDfN7DMdBqZTIWP16pcyvHto
0LPyOGt95qpXPrac166NR+K22JERcbaSRL4LpwxAC6zxSNdF4fmT4CX6GwHLTfgaQlyPbv2Gyc0C
eHcqYRzfXlsO9DsaOpFgR8FSI56oqHEQhv4/4gP0tlqkLX9JKzlakzxf0fAdeOTi+9uIEPqAKJMJ
Um+bNrNX52q9fFjQjHZ5JvDAUj8ZGYjtO5YNSTXbRl+znsjbu7+ruHx/u/bwWYyN/OVrWlpSge8E
Ht4R8tPu/8VLY3HX1gHHrpURWI0PTRFleDKQzNXlf3AmYa/BwQEttgwQPJhjlV0iZb1chdKrO56U
6u5CUx6EEvHi+YII8pTtZhf0dbgIpqm4vIlwESeFtRMfVmOsnS6iOuAwe8jzmbTtrGZJRirJNrvC
9i+Ey4B59DIY2p1Zgh58zF0wd7GHHXkhzs6wUICEdfmMvE9PKEYcMkgYdcD8u3+2SmV8/T9cHlBu
IoEKEmVG69pwEj2XSeSOktM6HuDR+XvC7Jw6it+gz3WVehaNa2rnhI2/iwQ9z+/OojXuuSkXdD1S
N7bNCn/2mZyNApX5zijjYFEXf8iLx0qN3sw7MZP/T9e3mieKdGab3fdphLEOgQz7z7WEq6nktcSE
0oEYkF+YkaF+lAg+HwICNwkj46KD3tV51RGYCQU49i7ns+/a0QyPTQHfjlzi6Z7BDNE8pvUejGyR
/xKRBJk/AkxwycCL/bVnRBRdoK21i2g42v9haYPrTvv1FIUxqD+BoGpacbzz7/yqh9j+RyJ6ryYQ
QIysDaL6NOwRlUNceWlWCUAbz2tMl7OFrex1gDHiimRje+QkCuvYZM4UmKGcMk6tl2QN+AhOMbPA
4sP0+jjKtIM0y//4tQN+cFpVboNuyvxWVEeoh+IXXDhxpwuSawtvgpaK9o/+6vAnKAgyaLL15ImQ
/9fj9oZCf5B1oI2sloaWad0s+6wy9OYMW3DK/xVQyvb1aR1cA8hW0hZKhIzruRHXBprPU+9/No3u
fg9HxTLYP9+ED0tRk9SY47wm4WctRl+91GbVGk+6IaWyytBCeuTYTsDVMsh+ei3XUFr9sr250p8m
Y1N/2UWvAdhlCLG4f6Oj4BWET5hk//Xw4UP1eYHUWsmTJTCyKfcVx0SOevs5VteG15FyC4yfDp3g
kcXucASUSI7metOGmmbpfa0hZ3s+zcbTWckBrQJHy3Rj+JFpXJvAlMHY0M2jHNw1zhq07GWBNdTN
ZBXseK534kl8mtzWjilOS/NFt5DI7z8St4W6sydfhmktGQRKepMHg3AmHTPxKJfpB+7Si4AxFPLf
a3LK5SgLjEwXIlN6dkaUbPZsuyD4SKBxG0NXaFZs0hSCzFxMZPQ/Q7IS9amOieh1sQ/o1s5RcRPX
l+JwivTBQxyCTUrZxfDGPRBrWSCGz4R5JAQSSvvHc1/ZqyCeODxhvW/gip8n9XK8ysQV2nEPIELY
scpwQnRXAcHoRzZDiOvThlk4TS74mQfqWCIpTUwFU/5C1g+Syab/nd8/hJA/aThLmJs5VZcjkK3S
BTCevXx3I3vdIMz5po4NwJOQ7gnSLo5GNb4q6qeA6OJ100qfVhi4fH6/c8FVCxXU7sIORUXn0W/Q
y/68Tu8qBU5yExbr2Jls60RrsKZWysaMn/3V6xGxIKpXBUBsTgvCzFnkk7QhJ5pFS5VO89MIAVrS
P3ajTYCR2zSRQtv8LWVCML0WwoPIP4pBC7ioh4dJKHfF2n+RDVwtaxkw4nRfdiO5d21Crm+ReKSS
U61cCJmFouMfvYPi5FtMaPKRdMoplEV2S21sl6SrAPG0h7X6utOuY0JLHaSAqBFiS7S02Q5iP/a7
gY04vGM4J+C/zq11iUZGMpJ4gurTga5Gjr+Bq68igimzTIsHLiG1Svk8yRVCT1v9jKuk29oKC+NC
FrOGJjsyEyjejesdir8sLzV39YPXRiKxkhCAVfz8EQCDWUSxxMsnbblsJxZU2SC6VKIfqh3Qe9vU
9IJdEX3RsklXAArG/yHtf4zuX7zY2SEpg8LFsbT+rJtkbZfXm5/oLdlBUBhkMLeuQ/11B7zOvlE0
X+V15LGEhEV3W/xnsjp9HsqWbTGdSpOnjtBv1oQrBBUmlRg59cpDjZJ7CwYpZc3n25b23bBg962+
QX0xK9Ol0UG3mPZUiLmOnf1oxQ7p+Pl1qY15fGU2SVOe0lAavERmWpK/dQF0+s9sKDW3N+BX+OQu
OguVnJDGzAbYRuVQ+Yv9ALP3NSUGT3/ypxMMOy0SYChjGxMVTB19Wm8Lxvdq0mgwyyjOH5zS96RN
JGSLE97F/h9VR6xT7A162cwE6OQBSS3hFxd3Dgb6bBy3rlnscs1kkzAERT3J9SWZFz2meTwKWasa
j6mzH6b2bBv2gHvfCqsPlN6LexbMyu5L+iFmaKr6UbkhWECydNQeCzuefUsnv4ZH3/aTvxNMcENs
qLX0JKd5RYu71qYUkY6qa4aV9P00zSmcGM0deg22Cmbm9zWtasIBFh02BtrOzuK5Tm8GbZ0gEGVJ
d4xs7kO6f//IuTHTNRoQdLTkXJKqKk9nDfCUfxElZriV4cdAGsZqEu6CZBHHWlyXkxdXwpnZzAwy
2aT6eRh2QwWYCyLfNJo4U8KfBe5+cs38N8bo2VXAP8hMdgfpHK/RqPA0YaBNLgz1vzTtjnMQpx8J
joonSlXlWGk96R0NQCf6xwctwVSuZf70q+wzbcn+3jQw+m3CfXDlcwyfCA2RjqqkJj4vWOohM0OC
bEvmveBrxprHe995X6erVcgjk+qp+l10jt62NSUwCL5P91csmBmYIz50N4mc2N5e6iYFXvEEUgA0
QpxjtICQPhZU6qKG6M0NyvjmkEXTXvYuUPa66MFAGAtR3uReT/VTJyHgIRyW7B/0mY6KeSwEMUk6
/lCWQdYLI52TVIqPOrf+tjhETfnWgVwPlKQmcfRao7P5k1VsxeNzWcsdUA0I4VzrxKMEwrjUJo0k
WfYsZAX8jvKGfK1CdxHX8OWSbttn+G6QkIb3Iyh89avVrvQun4U3FUF8RpcR3UWBuzW+Mg9tV41z
wpcqhbQq/vOWGVHR9yNK4M8ltZzb92A8oxskxOCaXuO8HcP5Ex5cM1LV2Mxt+GnKJue1woLcoPyp
EuMIo9c3RKuelJDzRFdqU38dtjnoj3mT6/ZmCSVmhQn7UH2PF2No423J4nwzFbkhSivEhfLFrmCD
BKj65F2hmRWhOlStEzQxixvp/Ud3YRAGgWi0Db5/WJWjDQFpt3TvrdPkWvpUc6L45dX5CEEvpo6o
Vd8mc1D06aHtB0CVEFNLo9mTIBfnpxroZmEtK6xzOZxAPKEzfSj/fwMUZaNQ/iz3coeuJ618Om8j
wTaKwlo8wVgWlkLQO4AZPOGNOgaLa/NiFP/gHUf/SicfGP498agZH50FkSA8TvryWiseKwjrWQGC
N0KlKnGujRJNDQLS0HkeuR5ucSFjLR8f3Vid4WN3IWEgBjTF8EvAH1gx8XKwBZ5nuNazIcezggvf
OvNVDOfEEREmygkl7sSWYJEXa9I4qfE9psGC/OHZXS8VHlPitlwm7CoGpFNu+Hh/FSoFkHQc5acK
7VB7AZuHxOdXL0/AEl49wu6xfBZRudQKHoa5Rwxzpy03j8OprCxISEDzkUZq/Lzepvd9VtOznmgv
ORAvJFxeDvI1boDDeWB7pgpGnyIglx+HKc6/iBr5B2mfYbCQjYVEENBOiM5PyZBXtc7csCHDZ4u5
3lUznaMRYx8VPe/skBrWsgjLwDd3Kf9wW3qI3tm/PpMfkNqdbVNYIo1nVO5tLD4G9IhaSWiWLG2M
BvXIpD4P90LCwKXm/S+DkMUoYKe+U9HMi6OU88VT1Dqog0CIaEtEYKsN/njWSztBe4jalY4jMtI5
8uBOS1k9HVvO5a3OdQku9L4cyETZBe+wtjH/EgvuNTh2dGCUwIDsprQWdoDGpA3GI3xKHRjYQjUp
ZLg61iix5VuaP6EhywrSk8gSsDIBUPiu1KaJAzmTWB5+HcHqgquUG8hCIIFclhQLoJfg2xFxa8vh
SBVjtz2Oyf4TroswpxAW+7GS2OndFTArAkSRzi0Myp7RcaDOcE79ZtC9LCR1gQ/PTftXK2Js2d4D
j3JOdGnVxqBm7+S53YEgyk4KlGBfqj6hgRMDreXY0pUIgslSpCChgqy63krC0jGyKfYEs9JlTg3B
tRVPrk9k90Y3DsIEn2Ojy+rYyyEoANol/ZlXPQUJKYch+94vdcye2+OoWhUrKByzzVc7Y7E2g6vS
HtOzOtcyEnV7GwrE83Tqy34V/yCk5cxcv1pDgJljTLJPbt7/1rKH/b9t+wo+ZR7QbsxUpst7ol2T
AgrfSnYm6UngVdfTH9sgCVQk78A4F50y79GwzDLpu7pkZfuT1N5lvzvKdKbDM0ex+WdmBRl7JKgm
r1OrBNRzoZdFB8W9+OivD+r+VuNIYfP1M9pzs0GreAWBuTB6NTnEhC4OiGdUS7ADaBLVrbltM1Hi
p0C4l7VfVRM9p09ZIgzUHArhjMzcs+lQU8gH+ZqAVmGVDpS7QxkB/CShbw7gwUDfSgUA5v/noJmW
uxW2VwDmp6cD+aVLdLqqmHxyJGkw3R6h8zpftho/L8PCfkbi+7BpTXFfwbaJhyi+U5Xp0j66ocL1
Zc+rxgg+hvS2dQQvgXiAHAIvU0vK1b5cKW5LxLR2QZkOf3FeGEpRrj/a0tIYNyKHb9D5Xuw9wzYN
6K8vjL16toX/hDv2G6a5LfkhEDAxnaECux/44/wH+sEz0d0w5YFGP9LB1zRdSd6OabPcmsSXi1IY
ROavOQfLG9E0T4b0WQE5dHSvlu0E0WwQVKgZ3zd+4WF3SrWChcYMCbKLhiT6qDyCOvLWbFNuVNqr
SI660/2p6ekijgEOWRz4APvK88KGgJXfZl8AgSj1fFUaIRrXhxWrNIoDWLBPV/xIo39X3D4y7Cvy
SuPhTam99kRcJ1tr4cAHsi0/Cx/JWyBmNaXlZs+xke/TLs5hv96zq/5osxPcbo5pDXVKBGqGKkVB
kg+5d/OZnqzVw4MCij5EzOW+ItIvwnPPBv/EEoCv8IG2LvQH7sAfJCvtTV2mz3SvcE8vtNy2riVU
mAjfrA2y68Dig4mTWbmSUH6KENpY/kItfCZnjc6H3ZFf6tkzpbaNw7HsHjFfz+IH4qfW/Av+6gda
6K8IdgSEt39KuRdY73TFccLGpC2rX4NssVmWlhwhtOMJmkpze2OAr9VI9vcZbQOlcmrG3JlS0Sfd
a5fldh91eVM/FrXers4dUeMLEqQRn3bCSmWrqpxnXZeX3p26L+0SkXO2LpRFlHC1hqxtUTcM8QgO
we0vmIZpI7ibXFLt/WRp7mONedLE8s2wyJYoLt/FXNVZzlS83aayV3OV8qMiAEuHGpBxXBxXQXJU
CJKqoo3t9EnR5kcHEXj/RdoDMy/obIq8nB3oE4XZ5mcEgTLhm+iQ8GmudEMYw5DZULCqHBIs1y0G
xQpAzKODLYj0dqVVC7XFEXd4AzqdeeW295cNCPGj6eOuRM2ejNcK1M1RXyZg4l5LgetTPBdOjK5Q
1QyoTDf7EgQbeQIxkJEmcxOzuce1CuKt0DV+MsnH98lHoh3wCXCPJYiVvW8b107eE2RlHkj5BgSe
1MPU4BXu4Fx31SCv6GLBFmy+ldJbI9MW0ujj6IaJwole6p5FgBoTyfeKleHw54+7VpIPlmODB3AJ
srrK0ivSeGKz0rv02qhRFOKU7hEKNxbTLnvaY9VzKSJj63XH9nOjatwCPh6o55/eI2oLt9R8op4w
kMPo3EN7dRmhDnXnKL2ud+1GGOY1WOXeuhJGa8+maAV6QnTe3pnMM+y6He+9+LX21uUIP/olAmpK
FDnp4CYibeQT1W4zqZP49aC5k9oY4HUw7HyAimPQNbHEqqNdgSLUL0Gb3CiC0Erc4spYetmjlBuz
PygU3fgPjO2fEnTiEhSPj00UC1v6UdpkRrs5Y9l4XyiHBq3pc4vDDtSxVgg8nRYHBQXjlAbwLfHF
Dgt72xFAUKbSLUZEK8KBqygxtoembyTBXCA2jQjaRd9FeHr6TbX7QRCawOQwuqVlsYD6u0msYcIw
8RgwhuKoa+KrcxKDbo80Pk8HiZcnZsEJCOvdoaH9Lfm5c0kzALpQkGljmlSSMkMXn1EsUKWBjlm3
rjsa4wgOnSw3n5pEBO2meDSnY7vNsO3a9zH57o7e/tnrJreyQFjqT64+z51FvjS3jTmnRf/uGLAe
Ygh8o199r+Z1RFuuA6yGCGb/98cv7BPpL+wGl65tlZ7VRbyCLwFmRbdYcTc00Uo0LLhPGdcbP5A3
TXBrapp1MRnuKHSBdBFpx86wuffkeWW0QVUWvOTbDTX0Cf81yowsnxL7vfol+JEiOVxJC7pLGlTf
YEkdMKty+4xAxJ7HTY1vU+mY87mISM0f2EeW45zEamDYvdauqaghIh8YubKHpRARE3iW0I6YVtXD
naam3x3lJ7A/R67aIzDK1if/dl7EX5K93GLmdLqSzPBNbZzgSYpr/jAeBo+bT0drnXZ84b3Dc4sQ
oY3NGMsh6+f9Pr0W3uAJrWm39iXrakuEo/gZ6JKM/EPvNAE7vx3SBHo7lCf+4guhkIC7obSEBFbm
vcZIquIB2bTBk0uWaflNS8utB8e1M4iSyq3ThQyihRRqxOoIncDZZQwnUqFwgd8jdGm2pMbPUoZY
E4DOv3/ZahHQh5pW6itfMbI8fDyZOtIYl/3fzPH2iInCb9DoEna2pZFW0cf1ViO5xo69Rph3UAAH
b3qLFR6txHTJX2Na8gCm/NAeqiH/rUGa2mG1tBfXt3bOGX71EwNX0WKTYmKE4aMbgVWWTFq5799m
V3WdsaSMto0V84AxeXIadElFTyUZLW4L6gNMK+GLIXDbkbfdCQJUVyBow+kTaB3faFkyZWAzxWrJ
jYUrtMJyZTu5Qx6n+Ge6Bkj+pmIIy65vSXX31/KkKY318QUuGQ3zel6orSnqSRxYIGrLU0xrlW8U
W85EXzJdJ+JKIr9Sjx6kLAJb6y39k9gqYOqGo0PWejNNa2DdcKJkiq1Po8BK1lTLTb066iQS2Urv
hZFXZdRqc1Jo/LsLkqBcuTmEXetgtuTy2MsQbRH4o/pIqzWfkvumPKySa3kGbHLWEQBm+sOac3wd
iIjgwbAH5QVo+uAbCHMJsjjVlL9NYFx7LUwrNZ/OfpGxAhPpwtC0UA7RDgF/fGj5loEf/uT6tnxU
ibFRW/AucKHVlX85DeT9wtlaMFxN99GeDF7mVd0UBA4VmAXkoZPMc+yYCFhaz5V/foUMJmALecdJ
z5cuprGtrmWMF5IeEoIo9yQKmRcnnGaILokcMJfukGZQFpJAqX5IwxhboL/QPTJvN9yYl2VC1z5S
v89+kxTDN1xZ9LfFcYJq+q6mcXdhmLUWfOsP37nIsvByN6Qs+mqvOF1Xz5S9MbkiuuMBPZn7rhms
AzpwoJ93JA3NW37GQtTj6IgHN0kxlV+HY1pjFw31W1wgO4JPlWQoIZkmSTWabsrRu02X0JX+5jXA
FCaWOT5GHyc3F3FnT7J4BCfjUYp9WYirwsiwZXKWX8ayehVgfTqoaxzEUKbN4D1WEUyrY0hrq/Jf
WwB7LH2EExtcsbe49R7ka8LmmbkhnG9Zat4NwMRUXkTiShpU0S6uf7LBLACs9cKv1pLfIbka8/zC
bE/iavkZxQSCjKWAbk3DTAsuv1u5GEWGntKMRUG3et3vWvRTJtzCD7KFqNLm/a7FqgMM3U1Y7SCe
IxJ4+DWp0Kn/96zOT8GyyafoaEfyI0fZG1Ibyz69DIu4wKAqCPqg8E3KvXeGF8jiPdR1Z1ZxPsGA
jBWJQ0kAIKWmVLRbwTjNtT+hXJQjAvx+BXsJtOd69Lw3yDnePajV9Lcp8uKBHhMJB6qg+J+SzP6F
1Iq/3X+O8/tDDge/EElDJWTaNthyQ89grKz8eQb31qunacbR03s9RGpAttDjgV/0uwWBdCIEflkj
1YCjyD5S/53zNPuwS2eu5zTvhb6C6ioKi9mJExUWyCzc14LYjIDoFbfVrsv279Si+EajUchCAhtf
gGDp2TDv+m8jXasY0NOZR/iummRDJcnsSQJGSHYL1EAW3UOc0ZcPwHwnF5wcKZ9dM1/yhKKxamQ1
4FXk7FUzA6fSyJJBImXqevyvRBOcN0Z4HAq2mftPn+q9nnsPcAD0Lf7uyfSYdNC/a80SFTJJQUOR
UGB5oWYBtsIHpAtHk3oPvJlOcfzl4Mw/o/a2WIZyDkPS1RSitny9FTIks8plvQFcIrpqbTFYfO93
0/bxk7JG3C8W1iLS2K6lhmQ2Lji4fvSLq202SusfTLMJ13BVFgegJPJlQ3LRutNTYO4Xmi8Joykz
nPDDM2jLuY/8qfjbucH2oLCq5vdedwl3+d9eX237bmWQsOQlNhLoS8tOjmrf3iqrecQAbmcMXtXW
cQDYBliKSNRK5EHDzI5/zgMKVN1wIvyv1sQZ3ymOQM/KwoXyKK8GbsGzsbdvLBh5NRMJNbtSjrCU
X5XlZrg1sWtt6rBUUZtEo1M6ypNlvndcNuIqHeqDPzchQeiZnMd7uoyDSJ/RLb/KMnelsTZQeV0g
ahycF9t3r6lBzxPXIKiwkw1SBiW1JjieyRWotR1m7MwRztkuyhHQ7U6+kvSy9kUsQfGvXCFGv0mg
h4wV6y+MHU7gDiA1ZGpGD9h8Sq2S7Gd9n7bTL6M/xgQqoON9Ct5ccykBN4AM1vM/2WHmlGSZqYNv
w7uFHNOZD/Tk2w6RrQ7bveNFsDUivrF6leRvf4tM1Wc6NZv1I97MBUy76+RXULBj1f1iR6UBZsnu
dXKl5qeRzeKbUwQ7WU2oixUus+oGf+TZaMfQ4EWzQVfnsf/nMeRtMk7/wAtOAgc3lK9lulNN8Zju
DrHUbeYEP8D8ZePanPIv2RAuI3Lw5do52scENoHkwtAuaAKew7G6a0sbAbiJYR49/qpnDlcbLCOv
VyAHhuYqTcyMM9pBXbo1Uulw7lPFi/K1KlUNhV6tLTS6W4vxImTxbTIAJTBnIKsMbM5JZHSrt+BH
aaSEIVYK84hiEbjOtVjGW4c9cElDPgFDRoFX6R2cr/SDtMEAXewmJpF6M25dL4WAUDfOkRtmaxKr
1c/AsmHYIjYgCts9hQyDcMy2nTH20wxXFNbWsMOwFFL2hn0Bn5s8o376XFBUuidq12Hn7E4OQpdL
kA8zeWnjKv2FbVnWkyqby9m4GslcvbBDsDHlX4dsmJei5KUPasldB5CMd1MoGIr/yk1Yuk13rrKg
d88ehNj5k++6iVTI7E9LrwqhwXfX+IYM0j+yq+8DHWbcSismAvdc54gwhDXLHV5X9gtTOHlzYA7O
Tsd2/CIS0Ng+XeFsBOnpYxVfEtbZLzm3P9WHt2CMpA/L1PXqVrD8Ot4jf/6b65e0Kajez5hwcl0q
SgDmzwyq2xiVMDAV/TgAQ9rKSsIytM+IINQbRSdncByKkUsqHU2A2Dy3ZAo6xuPXFWJmPKqGGgvd
LBWNzed+0IUfO/U/ownFLwnAi2KgI0abqq/amr6T04L9iqyQEfBjkpwqfLV1FrTljQL+Qw1BGfl/
xf3SM/eeP/0MMRBiqjU95SUMRYgxr5z2nyUtzoENycPpXpiMhajH0lixThQnpgmdBQj+DAHR+KYO
8CRf8aurX3+TK+xc8GR0o8s7npn5eypcVTQkrqsXaayL2kwtpk4c+eTl0/4azej04RFhhkIsACop
dioDEfCP7HIDSr+Y1cux8bHj8FIoW3So62QzD9D1Na0LHaUY/USbvGYoarUA9CDSt2FzX0MpjgT9
6FvOgMvspz7Lf08swqoCpPfmFEpBbsJTNmsuXwjqR3HoHEteWh5UPZIlT9XDqpW/TnlHyGoUmRko
wJ1LMbTVsEkE3Wv+VdP8lf4RehElfpsQSDPQejHHGgI9GPuHDMwX/r847J7mAopm1cemVnVe0Hik
Jf8dnT28pkAfV6pbsJ9KcnpIJisjq9AjDrhXPPgJuBt1fNjBLDZ5VykBGTd9Bc9FriMHmAeTGZcL
MzzIjy32HcKhtEuUsGkHazaijG/XQPNO5R8eXTV1AC3egDe1skaJgSzqpHYgOT1FmXtyXWKer9g7
+k73P9IvqJq7nJqdwIvM4e/QEfd0ncv0ukeaT0zv9EA0pT9DEBvkblIwFlBXWUljYlzZVopADiVV
+VAQsQdIVF9ruBGzZ2t9zzgW69OQbZr7E68V5dd+e3rwwNWNqWZIO6guMyboKIzsIYxDox5okeqY
yRhk+THYiqYiEsBhBaa8gpGxV/3uFXwlVkUc7n01BTtVcNddL9xAzcOSJZZiCUDARuTsiowrARnY
QhQh9CsYFxo5l/UN5VnzilDrVBj5XFmrAXdrOaEShCrfiO6DA8jKeyxA+kJVxqBU1AqUiFvmTTRP
swglfiKoylSwDmE2tEMJ6v3/pQL+6bpob8C4WsOJJulm6JwdN24toEnkeVaSs2hhB8uW2ncRho/Q
8lm56qCVlVMix3+Ajbloalvo8aFcBz8TW04aLZLWB0ayvIn3VavAnTGBerBgjW1HAowol7uMs3db
0GmC9H/lImgYPd6v+OY0cSu5YUs9kbc+it7GAml8/cN/8fOYKmdpJOiX9+uDt/0DZQ3I64ns0MkF
JLLJpcTCdrLvy4L/0SAoBdRvrC+moU8ZGtamdBEq6rm3E7pldyn0vD6Rig4uJdGSAbhroUo0f/jy
SIhUlUabov6f9UrxqH4GfHoBQA4rY0BNq10LteQampAjMWTgbvIUu69jwNQ7Lh8M7TjnMhZAVgsp
UJKv4NBbBW78Xb/F+MwdQQsjb6KCPNzPASefCrKfm33cV8X1Cu7JuDi3+Oo/U8wqnMKkf7CRteRj
eQnxVRktHMCA+vsk22ZjbhotfUvvlyMAy3egwViEwVHvth/ErcEsaUkroTWs8QGOrnXWOAOxa6JK
KivaCJglGOAvEpRv6UMh1V0PLSVHYZ8CgUNLD4S3msMDLpEILADeycG7rw0f33h6oBlhw+nOezm1
O32YUgJqs6t1Ng/H8deYTFBzFKbPn+147vGizQeQHMcF5endsLq4eznV5eP6tKFimmT2VyBxCwTJ
6UBzI9OGT9ksW0fUU/P4Ol8xsY6KJ16xZJnDSjQYXyBma0tNm9t5K6UcraZazKg7dRU7GNzqE7Ze
ryOC9YQ+T0w19eTnERwwDacRS0LBvLBHiuZGP1qTgomUufY4da8zdkGpUUSQ13lB99D2WSqeP4Wj
oTv5F2i1UH9Xry2gD5HCuNqUAw0qsD08wh3qHeT7FRNnL8CZZDPzuuRfRtPWPAravMSTRRoWevnq
poBUnMLdDA+F10nvKRIFpCn/J6NS+V7zGexLyQunprOkFIf8JbCbSXyji/3VAPo7gLyBGOK6CEb8
w5CHS4+tRMQFmgtNEKc9Cpmq9B4R2vl5lc9x1w85KWovMmmUP86YvHh/o5vSS0bgTLH2x9ULDheH
upxV+3BaT2H7ujkk0wCkmxPzQyXHR9mvr74b2P00gCMvlAJtGM2iAMH2+2sua9k0YjyBP+5bYr1F
3GYEZDtZ78oFkAMnmzBJqWgwP1EMBHizTj8WsXysFHj8eS3/3KcaZwx/3eWDC4BTW7UbmF1szGlM
WsntkAVihoIr3yqZ4kllskX0ueRYyhC8rfiB44t5qBQN3KIUb5M/51+v3fMsdUqEpnOk8a+XWba2
XA3SumeTiK7tfKA7U8mhWhz6Wieb8HnUIaHsrYNDx+LCYlm98+C7mLEBf/zG0xyVFjtQ/9igoYc7
ZYt3a/rZqxCNtkWj0Ze0G14ZTEhmYMm1Ve/9lkfsy5tS/ro/EYAV0Zn2lehEvohi1fW/WYHoXFl4
CMTWferb5MZjhTIk5XZwe2jIGO+8PmoRbuFMGhq8G3JeK6D1edVfmy9p/ZtJOCZKFRdSxf4X31el
3WP1fKyc5OBnHIHCJggaW74NKmRPH+K2iAbwQqSFZNx9QNO0ErT2iTDwrqhrafb93LCLZb0kE6M2
lhl2jRzpTMkWy2vxghC2pisxYUyE+bMa8tD/URZRtdTrjBt5KlrK+RiOSCm+dey1jRjmngypzP8D
zZ/WxKF95WUJzGgRXR3sWUe+jSOjJbP8MEy+qjASWbzaLORLLiwQ1rG00DRsQokSodBEdqoFmKxx
i6XTQ6VVnMGXntZvews4F0JfdsUJGilQvZeOjf5wZHh24O2cIidgR5DNL9/Oio3rTO3R5nC0IBnt
SmJ8NeNAa3B2xYxGcl+XyS7rPoswd6uR2/u056kN1XYzLm81ZeOTNgsVoVt9T8+q1/kVlbcw4Wzh
SA+3HZLyUisJ/mQgeXIPTFSYNdWk1A9vrw+Ip44Zv9Jjl2hkr+IkfO6/pPpjUq2IofNZDnHj8Hb+
rqlgPvbnX7+uOeA4cV4oTyAGngPg7FlQxl0PHRz2i+sor+jfH+Ijv0Ul8ySQ3BII+gVUK3sA7btk
LmVZZ1ddVUP6kOGDX6Ncli948kHF41VJcJgLyx/4Pni/KoMuqEZGutobxLgmQBhuNjDbvpP9YWo8
kkzz+dvojJT9m7bMJutJT8PdSuUbz70WUrUcIKZLrGAFrrE9JyfwmkqQ4ZinpM8lrifpZFh28lRA
Zf3xa26ZoS0mnwDOxQ4HBfcGCNHUpUtgotd/THV8a7zvfoUlXjxkvwqYNoy+YBT5HEAuJTy3q7k/
ksQHu69QIRILU4xvJbClKbLg/YCvJto+cu2J3oY3NyQh0wBKESm2zPTLFCA0wJiq6LISR0Cv/nGD
7mWQ2uMxWoyjJD+e7XFkFNSHzw06XquHfcCZVfbjI3Noc3vs67nCK9xFTLozBTs/2L3ZOLF70xa5
aMitVmX7S4alRBz6GtTADNhMdGMrpORe7Jsq9j3RluOKAQzal3FsrOJIi9TzJycPEqGZNANQqium
YxFEzJ4tfRio9S4FsG1iJwSgqCYmGtrVnPwicy8reichPMJGL1GZV4x+EGrHUJsMs2pY9ygGxJMo
ls0oGOpaLgGqAiHZnm/kw1z5B3g1RbdVgyFnwVuvFT/1Qy0s9toZ+lTxJ751s7ZSP11YbB0d2Kqk
JIJA8h/NK1ld1uDY1iOk7jqoY5vjnIS8SELGZxocMZAAItuDsMJe24k0aUNWGKVF8r+h+ITP0mba
T5bfY3CSfFM78uxu0DmGltXYj1l1ws7LhRoIWhnlsaR1TbNRR0wSCTk3izD+VJzG0IOliWT7+fFu
Y03OnCS1fBv9ChH97quCG4KK2tDHGFhok16ETHoH11PJEItyqQ8qO3aIDt+Xagn4MLUG7URml37F
rh2MIbVIpDF42/DA+xxu9yXqhuZsaVNE6Y4nnma/JClm/XMeBqK6qsQ/L1okEAGP218P0Mm4Fcs+
fydmeivcA3km3vbiWnYxb6z8I0CN0z/uuU+TAsDMkw+PeJ1reFw9j1fwtI33yf9ix+aUdhWF3WbY
64NLo9c7ht+i6yBFPc74Q/M4VHy0GrDdB0NvhgMHlT5/LBuMWhV1QfJO/nCH9jO1DF5TnPKWI5eZ
HwkrKWAt/Bxw5oCXv0rndYK/MoZW7NnTMtesvNvxskUfI+7P0+L6HzuzycNdLeLAmKX8WiN96TLS
5DR1slOQW8vLAbhRE7zRpEPN+eIzpO+rpSl7TKc1Ew+nvYvlMICwAuMiI7QD+rYmdle350hNXuKa
jSkWXmThiR4I9mRSbLWDt0T6q9y2l1pdqLcdbvi1gPrv9n49NOMvcIPetK9axvdMcKqfOqaU1IPH
ttUcP5PA6qEwr9SwmwaC1+Q3VHwI35Wn3sn7JDhX787FwT1P3i2qVunuF6FhD+JNRd4YsP7aBZDe
zfchtbZxqar/u5RRFOgps7G2tMXRKEh/8seYsVGX6AMybBEPHIIhUxiy7cHbDIsi3i75RHGXcTRG
w6x7NMVXi2SYpMTyic4NAxRTh7aOmytBOxhXCYIberVjfq/6s7R+aH9XTBEt6PNljuX8Lhmp+s0K
lZXNwLYvw184ISKdG52rN67t9ppwoya1P7KyKfC1IUirAdLD8HyBifimKzZ4JqcgoA08tPnHIuwj
01NHD6AoyuzjAtAXcPR4c62dOH8HbX6oDZm+arfo/Lz5cccJ06Py9Z/wKwfAvw4+T7qH3qF15/iD
MKNqQzvH5YffSE5bdmlf5/j4RXGwoBNDHRkEs6f1Of+vqCOGkWy75ghY7LZnqNm28JSC7i//TGi0
Y4+zzx4Eh5O1RkewHUfqvr8BN91gB3trVIBlsDIqbMNv9OfuiaNEV6aZIJsb9arfoLC3SbwEUxEh
RDgMS9Tpdz1qMW/FHHpR8gThGV/Cwg2rldygmaToznkTvJGAPG9WLKHKFKCXCtawWRzR1nJz/xCf
FirFC0vHNfJlHJryh2f6XXM8BWLd9/nNfqKLSSEpUUQ3mVklhBsIrhTpHgM3zyX/bigldHPh8Ll1
nB4DoFGMwHymCQxlwlNrZHt1BJJiMNL3gTiuJWEQd841JIYlejcwmxU1c6QGXb37cXF76Mpm6T6u
euYkLV1gjLeIBZt66+CIAqjWAmj+KUcBoV3o0LeWOXraZC1rYw2+fql+QOn/o/KpM3QXono42zEq
7VA+ZBO8v40qA93BJBo+3KyTPozHcmwYdwFo2TF97TlCcGB3zz5CNKSHy/Msdp+856X077ZUbn2W
IWBDQSYpB9Pb8YfhBWgAEfxwAapru8xQg38wzidI4E8BFPqeCEaXLK3nKiaYqpHPEz3W54QT1/lv
JGce8NH7nBTJchMIN2UIZrCnM2PImFdarhIzW7ZHppCdqsCFXJd9AzKfti/ghOqtkOKyvoZ45dDx
W21YkxLn6wUCyx5VfYqEwlxLxN/L6qV8Cu/yRhfBxWInkVFZXVjlim3d9anT6IM5sgRRCGPScqR/
zGrb/9EqjStDMPKaevR4L06NqyU4g4alzLaZTcWoS4HOd7rNFwu1kSmOGAcTu4qECp6pHnb6CoMC
LcZhCeImWPDTybhypokiYllKRXoeCgaa4Mhzst9sbdDkGLTfvMoLbRUDdgUdglJcZjD4+DlAdR0d
o5i6fvIl1yUOh6Dxy9flhjCNZSi1I4bHJQzY/E/J6hdoRhh6ls88Dg6hkxBLEvLd+IqDdyRcpWfb
sPXXDmVrrSCUxdF90b+8YVfO0TJLoAqpBYJsqBiMnt5eDNc2/VQ0owyIzfdmj8f0iPGAN2H3/paX
eN9FDlvO+tevjBZVWu95YdmcQgMcZBP1BE9AJDePjeKtOF6agyO3AHt2GyFEBGmGhut+nyp43QBc
E+/Jdb1PrWqXSgbvzlBKLs6mjVO+QNUTJ+xC6I1fvxpPv1KF3Pyq60V/nsscy6w767NHnSylgfor
rkDKGIOeauMr9tbYQA1XASDCAOifC2vsnDz1rbB6a1QO+5mrUPlmxOnd5EbrwiXdx+Rrle0JpghK
tuN/y1UKCop8nDbVxumFb6YTvWRrUug8AQnEBxkMBiqJkOB0ZDExCrbBF3h3ZEYK2HqFUKUuUhpM
pRgM+pVoAXp3COEL0bVl04ESrqEJ2tBS7Wg2ruT5WFm8R00PILAGecCES3lb0OMrWQri3YBVsPvG
H/7AfN3IHPDVDgvXRLB6Vcv8TeMAVT2YzG8jBtpUHoc8E8NliW88nF64WYCbCXlNhelP7wXbPfBj
y6xw2vvCPF1pAMRrV21C7UemQCpM2twpVufObuQ32naOKZfHCXjxIKC2cs2dFGQGo7SBsJK8M7dr
IABzC1CPYAT7ruFdUPmRX7HZ04DNhbMbLOP831Elx8T00Gyh+2TUPZtQbR6gLiLmlImuEhNzhmyE
ViUTKN6q71hI7PEuMKV4jpephIf/5mUMj9bJWOw6GRNPKMEzPOcl9OgVkDWO1bc2rOY4CC57VOjq
fKIfIqZZik2KuXh4MW5IpovRzwzZOS/5Yoei1O/sfdsHcmVgIljTIUuUKkdRu7ylZoY3PwKiZWgQ
5WrlhmZ2mFlNs7nsUxMnsphLZWlS9yiCRQJmN0mLAwrWNYcKTEH4Q9u1JvwgkWdlL+b1QmNeO12q
2k3a8LRpkWMooAYMidSrHpn7xDtc0uwE8YsnogXVOSwvPCKQANWJ63ixm2J3mSMGVMaDtIru1STl
VgvaGLgwwsEw745XSHK5oNZFmJ2ZGmlOtnJO9xH5kozoQVPZVnH+wofFGpGaz7lgXVceXCpkgscI
xvrnZmlR2jUmIlJy2vUZGVvqyDjzZ81oTS/u8/JlTT9YjL6eAPbgmPJbtWC7HXpdqPFI6FljG8Hk
Lmr5J5EHmOtHxt7wf08Z4hSFUApQdBYh6NJhWd1slwqDyCz4FOoAtNZRe4TSkHiZVbhx144m9wms
wacAWtp7f7++5Xr3bKc1sC7BPVjwmgDrfIcel5wavzi7qQTV+LQcx/ubhsWXJCT0k8q+z//DewLu
9rxLJ17KJxsdoa5jXK6Iia5qUjIGxv39wGQTUKeOv13ov0GQ9h1YMm0/7j9KJvl+Phxk8rCfkEb1
QR99q/G+XjR3pGqkxUqZSOSYQGvvV1iGUbB92+IbCGL1EBhiUIZfV55a3l/vAVtwfSgwkSypRs8g
w5fdHDw0yamdIRYtX8WTZh+OgIvwm3XGJVBa15mR7+sjyKHN9qZ09WE3R54SugegAeG2+SPmxb/m
7eV9U4NEMzhpaTP+uu0vjS6NsVhM9f+vwo2vSljIdshtSByblixEAvHI2i1j2wUzOxlU6W2Zo5f6
RshrsgqhHWIYQ6i4s9j1rtfYO+bak2beOflhwO2sdtHjP50WggHHcy4ukz8FSCInfffa9bZZIcAL
IWnbjZyjr0N2uEUt4vdRk2K4uBMrFNTS/61l7ZBUyDp6yLlHpadyL+ZfgMmjy1WKB/sWxNkGt7tP
SxLTDnm77eTVI0uYjZWokyV4DUf0lLVgWk/trstnoISxJ31c84M9Os6REUwlTG+JTwk5SOGrFyzJ
DzF/kPp2L5S3ztSa6Q5OA8BgyqIxhnuJVTuoZ3kGYaDB+fjcvEPVCJnS6XYpwa+VD9J00P9tSxhD
k8o5+5fBtMTzmOUgtECc/VXSwlSVl1mvLPS14/mLgkZ5bteqd3IH5cWpPzge+qyUPTzUJTDtFI4H
8KkljIaWWOx5Zvz2yVTzvTAt09gn0lhT0BUIU3e0UBDmyZjfDr2q+yljV/InI4JAumklE8bZIDqU
j2LFWOIGJhhqGu5IyB2SalkmLZGgxWUvDFjzYyva0/Lu1vD8EGvY6hP3XY6JWaCTUaiT7IS66QDw
97+yqQT5FDaoVFXazYfh1WBiE8V/qdg0etlWTpK2oURLXjdEuMcqVgk0/peC+w2My9DKVmohAk4x
k31KcbvVXBafn5yPF01f0kWu9X5LKmd2ievjvwSkRG6WOr/THtaJ6HrBpuEwdlAzmXNqVHoBau/J
on1WW4zXJqiXAGZ4Ih3sjtA8xNoq/JdzjJVIdenlEEmRpv0ND3MT+6wWHiX6aTbxFPHM9PAKuXfY
YIueMPHxv5457nebhoYSUNWneizKFYeH/J6S6xcP2zEti8Lb/yOPpJOMcNa7sAB6b4tt9e6PyK7Z
/Blp2mLAWdDATmFA8wmViI9dN0af8bTXTMZLT9bpS59mIJHTNmZkkhOyf+NxfU1EUaENu2vRHgyE
mla1pgHk9bw/86f66C77FoyNSomLUKYGiX/Ft+l0Ez0zJweGSlcLxTGf9mLtD9SzPIUlQzGE9m37
s90BCPL4nQcOsrxQWfUVHo0uqAC5MQsyK3BNY37MI0WcPh3InE1filfqLQQOS/D37z52mSMev2kI
riejQkZqiuyR5A71Qks61SwipUHfG9OGLjXIc5/9M3WSEJNoyYkvy0z6kt5kjDliG8tNoRvKO4uj
qG+bMwLcMYWs42MACbhNUFXvFOekPQrh9GRTkgaM5efivs4nwEMUGz4sW5ocFixTsuMLQTSaC5yE
lDX2idCJNv0esygbykwuvw8M7cjNhARiW6OtvvVt+QEy8MnZgzEc+PwHh9hZNOwnC3y35hA38lci
wFspGOs5m2vveeThNVyKFScRmQSyoHvKmgFxm+8NnE6myYg/49mGd0fxfqTsxGvvlIhGgwmuH/UI
C106uNikVcdtlnrzjKJAYWt7DnK7+z4RLhL3XKRCTR1rDj7/pkZTM5NWnb8W5O2fLcUHZRwZ7wUR
VqqizyCZ7GMzIyXEHpzYkIPLID9wLOav41GbBE4Q6yJohqCeyokHBlwqjtyBArrFpyb8pEQ+1hEY
/c0wU5oYERmpdls0cx5Mw2WD3Pt/t0Vo/DKCawkqgt/aSPr4SUAiBlHN3eztP5nKw8/YL6cHsr6B
SYv8YC+UZ6mCMXDvLq0ULDZ4cmI6r0A+1gbZt1H7d0eKcebz91h5rvuc9sCvOa/XiSGWCiNZ7rBa
85w3TrBQd5mfTk0OVdAEYRbyfYrl7/NdHWyseucHl+wdBz/ob7ygTMr080eYNsqmmu+dRqcYS4WI
xG866qLFwwaf7paEzBgTfB7qhR/6ARFD65paPSvE23XBZVLpTP1Wf1eRDm9MLcDcwoV5qCokPbGo
H9aL3xmFWVgQRZpvqF9xMaowXcXrUncrD/oH5idqNdIgF/fujzPZIS+IyTxXIYMyV2JTK8lNcbmw
j4acPQ0TG1PjuExPNqudv0jSQgHUpAl7vKY72IPhqh/NExlDiqLMmAUXrwc8Wq5n+EZasOZoWl/k
WRkynGGSsL0dAdFvfwneJgSO6//3ovT+8ILjuXrV9xdr9to2dCfAZrHGQZjOHUAMZzetE7yPqmVI
6ugEXDJh77S8GoJlsM1ax6QCQXKYTKQsg9V9iYB6HgmbZwbPbs4EQg0MT8ackoUVJugpQYOmlnpE
ynp8amqTT+Tku2pq1iw4uhEnvVsfPQYefmtF2POma6EwU9ajM9pLOAsCI0xh6H+Zxotvl+9WENpS
IHzaXJhzIOAMC4CAFjKrk+crg0yfMQyNK6O7EJrKXJlTD2N5bpDwu6bkuYV557oFClrh31EWqZFx
QgkXR13wTAbF4+0CfBlS0T7BjBzJXiZ4H7o9Wl12RBy8z452h7R5zzUSR7Bl/y4y/A01Q/JRb54L
vSjX3d1iESMl7nLALzs9ZwR5cm0olvxGED0/5UAyrlnpykS6JASCu/tWwLxi4xsY3m73sSMWW4d8
hs96l0+lehT7wVjoMSnU2nnJ3jfX6Pb5RV+rbjLkD3iYYRYBe3fbPPXqWBGrhEdNKGBqfzlR78NY
rroAyUCTVM8RZPFxZks6KHcYOMeuL9IIvT8mjjYdYfh3AHp3IaNqS99MI6gs8d4mIsDR6k66b6R5
AH9UO7PbthP+vtWVK7J8BcTENogFV+ocvbpVgToZvXlDNdrxyVbYpuyaRVZmsDU7DZwUn35Ll3V/
4nmNQd1Strfl8laU8v6MAz2fLW7apzpmrF1w5bbPl4vThMa/q4lgvrZllkCfekD4cVaT97eX1dye
1wgzq0W8OJZGbJIEaaChc/1yODMprEhTeH8E0yxwVDQ8my4V7JN+6G6/xGJDO/N1r7DQKI1u/XMQ
ud2fjOisl7HgMn1Sw5Jb6+0nsIYv3d1HHVOdYqGbxNxiJbfulBKCDvu/YAFZbdqug5XmOrq/9qvJ
oPl1/3VlqzHWGp4RFMHlAoMiDXLGF4Iv9LlbzHlVRbgE2qZ82jSTIdWg3BNpdTMsWR60Jke7g1Fm
IIS7//U/zkaFL0t4pIhbzOB256f3fIPQiX0mmUFcqU/J7vYW0z/ImEl5o9IJc9HzC6AIuhSfUowH
aMMS6rkjbj93sTC9ilXVn2uxkaFpZ8ZKiDiO0Ur2t0EVU8QOVkxUcDf0i904Q1xlYFLpwe63Vpdx
1B2fKsb3+LuNF8Lc0cZobPCmVVHl9cn9yW1qyyjZNQsKak2CdaWFBN642+CPFtP4AloAwVXbFY9k
a0vNT5Eio9h+bl18rBi2yyzr5RTpGzNjW4nFrt8KOpW8x43ebK2UWdwyPAWXvfbwtVS/O2vhGkhN
mNBcd/OR1HR/slVtX3UXlmV6Q7b4EgJRPNXOZyl39PiNNX1pXeQI+s9HrtEgG5qMU1Iq0gun6v88
BtlOYkHNBug0pb6uOCMRCb9CyjUyfM6cReZqrc1+41HbYaloUTwwsJnCZA9nWUrRurD0ybJ4g12w
qSlcJ/Ias8pGsdnrRyRe274H/JK4O3wfQXujTw4+CravbUlYo74o2BCH7fWXKAgnTo1FHqN3CST8
bSNbSfG0hjG/9JoxD6IMgBw8Ax9xz34q1wGsAw1xrqiqwyzpZ0VoZcaZ33RAUaxrdydvcjmiyBj6
baBDFEBy+w4GSORrxfkcPNDefD2JrhBcuO7B+u5lGJWKtXqcwNasHPkvT99QfrCtKY9zZyahbBDo
470tr3vyl973HBxL32IFJEOE1qLqGITfn6epnXSbZhge+s6DH4bfqPXYguPYxXL2roAqhNeWEH+o
vVNfnRRhQfswKxcbzMNzssgQCfiKiVDJk1L7D5turNzSfBLOjFkbOtKb38dH/d6uqnPVULY2nKEj
hTkMtuY/Mzv0VBBdsbjDM4GkXiPUy+fHh6oxXrdJl8NG0v8AL1ekKISx8wAS6FaVk77zqf0X9bT4
sips1kCCwPghH/wQI90KVjn/2SIRGIvRPglGX4VmVuXuPcRedz1ojgPji86MdaEQ5vQ4x/LzSA3s
Vw1x5mUhQAcoV/5qhQ3ghUdwlWrQ2y6UnMXuVezagk7WEANAw3wEHyROVVEAChQ2O0KlALMUHO2p
BK+Y0PqVR9ZmOVpzOjU9N1VduYZPeIYL+zkevgntTz2fVgyIhpBvJTFuhgbJIePbfD8f1V0hYH5n
W7qs97qbrUZZOfYpD/RIBsB9M9frHksQeEB/sYF1bQoReOzJYcZVrLJiPLuSJ3C8As2CUXzppWSR
hOG6vu7Qx655Ixl0RsGclh8d9ULWmxkKikRwd0Uaa2GtMwBD1sJBiIV7hoeuEMv1wpWC4/N2o1mJ
AlgToUiBQLKXDxzIPfN7zfiFUDhUucPQYx5P1Dkb7E9WGELa84YS6OLHzpHyahnbCcgQzV+4GKWr
JFhSDgM2/b/2R/i5AZ6OICtAXEq6sYHqpP57uFPJ11XlAfijKc+jYEyW5WQLfxTunqCHfU5Sjay5
C9k2UvIFFJzz9hKXieK0IE50BknkxNFSq5WIXB5/R5KhzCPQvOJI36AY9ci14p61uK5lOPYGWx8h
5zQ3vRghNdvk4flLKPWUQlmzaxsJWmRGC81aISwjVYReceWkR50ivLyev0F+Lyy7U/vDWyDtTu/d
KZ0AbXjW2hW0n/qlyNaCBuc3csQt5Yhtv39mPjje7/ibTM4AgBk9YIlOdbf6SnZf160v7Uy6zZuI
WXwQR26myl7Upo/24ZkBI3NmUspDvt4VuP35BtBLj1UfYINK2yz9U/tftovR4HPATRoY5fHTw0/l
eqVu4v4mh+ZrFbSlbMmgie4dMgwX7QSqCb+YB8ZDSMHQvwJ4Tjz0sE67DO3PL08wVkVX2zlnJTUD
wjuUPMxWnqeYDgUkYf6rTh5tY3wn9cGNVWLMkQjjSkkLYd/ZsF3qhL/W63banp8JoGB8QxnZHmIK
R+w6nqV2mx+u/NDa8HkW946RPuC8pupWXb1D/emzb1aKilJ1uE0sk9CUTtvycOVPzFHGpi+ppKeM
0bUBadwGLQU85srCLtw1g/erPRlW5WKEZ6vf1PeJrjfcjqSd7L5iXv1zma7m1G0N++yAGckuuV84
qSCE/QlMUf890vQ+N+zc7twChh0ETx7bm/i3TtnSPpI19IkjRt0H2dx17Fo7bp7aBLlQzTbrINiX
Kvp8T1R/4VPROVV5hHGzqqa+fTS6Cr1hRL4+aMsTl8HbdHYGhP6am2wDz6AJrksXmoKH2Eg7dUci
WYtsHDrQ3AIc5LwbN5XBH029pcGY8qUZeQ6Z/5LmnNaA2VaaJxSfqmeXZzlo0tWehZXsYzkc1SXw
In5TaWtshN391AKEPSs9GYCJQTcVELRUMmfFzbm3v2n5IGevAoipw7Lp6QHRfkaEFDILdYO1SiGE
yqI05o9qRARkFyvmSiyNQxNEO7XwHBqTLp/D6SOooalmvJ2hU1/71LmPhs9DyO+HBTEHy/KJ9lib
AgZoNXzf/zy8Bst+bfG+uZrhGa+0OTJLmtdjd+cZjC1+V3PzHMmrhxs5oTtRqqtqwqbhLJyBrBcu
ukdxgCJIglmeP3AtFcs0+rT/xSWWBM3IYjBmAVDL0JtnYGBN2Myt8/t8kDwW0UfDfXGkZAcjB37w
VVatnfgqOM7YaS4Fko69Fq17C1un0IEmv4TiWsfvLQDUq/WAQQCN/BOoFsKOTUvrkEmKUj65g879
0YrqTaIYrYLe5S9YCwzl/ZTwahRZRCmpHvF7eD3ZgjFm3KSXJ/0QgoS+dOhKkjhYWSPYMfcsaanM
LWtfgoVVF9JJUh8QSGGbSYlDBvCf7LJ3yNkZ8PB29ibTBzimEPkDLrK6DNkddiT6XTvKVG4ykCS6
QisQfJOEpzzq/OBpNgdQONzWZ+LBujwLb2xupK5Rgw8YM4iWjV4zkUCodWiJ4iyE5M0MW6n04mCf
NXHHRz96f5ym6h2mzcAZLsLtJ/ovfVMuTV44q37qyaI+2ilXWBrkBINrxp1IrVsrOZu7VHIZbJGb
Pj5U1XD722/Y2Pva9p/whIE899gDbVybRoX3JgUTOjnI6IA5ZROaiMJYPmAvxFSFCyzywfv0DP2U
JOz/QR/SMACIEpXZiRuyUwAMAqHUqNtp+fqKwAB2h7aMxpBbg1lcSKiRKgdfAPZsRZByq0cyAovZ
vm0ktb3nI5tTjRHCvzML6aiaU+BgdVtwKMIO1gUua/zj732p4AKfdwaGA8gKL3pWlw2A3s9R+M63
61qZendySmBIs6r/E5tXn9hi23hERkiFW9LEq9/XvvZQSTc9Fz4yxm/1bRxRqZ4x541Yqm08mMwt
OFOIabug6dHNANscfifQKSNY5zFmVx2FirWJZfhY3PH1wzcl55LP4hqQnstC1KrW49E+gokeiIHB
nST2YdvX0w6rq7dHeZoaqsZqNsGaS0S0wGC8OwfgkI67Pp0t2spG+KmrOigSSEBHNORMZ+7ojqgm
KwWy2d8JHEJr+K/erJfXboEa+1EOTNxjkhxKIOL6aL2WVbksGt5sCsgv0JTCUaxOGbHzliGxGpf7
M2f0XFwg3zLiPjBQxJYLJbmwm1IWYl6Q0M04gBXzlE9p40q7nu0B1/fiNEDQ+u78qQBWLHh/5Dpu
V32i+olu222t3bquRPCEcMb6jssjT8iF6NDwPsXSDvVzdLj8uh7oKzPMYLguTL1j/SdB1NHVqGGd
YP/sFnDsDb4KQu2IFb+d8K18/2fQ3uy1A2U1Cq2LG87aZLztdmbiK4nl9NbknvZTEuknQqI7GBIt
yvEY9njzpuYTqImfT7fq51eoaXtFrF8dJKhoOMmVH4O+WHaYCPtbY+GN8EyUYMkmcwRPELaxCwLv
uZ9SKK1YYOz6855CFXu03BsqhsJ4Dim48znFIJES5Q4QGrKh4ZG0USqND9ys8lUgl0c+N36/XwU2
gTb+9GQYViCAZ4z2Ap1uPZiNd4SEH7lU9JimjrWoJFnmSjr+KXJy7vSKFrFXDYD4vI/Selt+PE+H
8VLA5/ncHo7Lpfakub60RyuFziDDl2UTc7HNXfILwu8Ndw+18e39Au7GqkplCHP8q+HlgNPZjD1O
SMDhX4mtpBWzz0mrIKM4tv3QmWxu2Wh+NUrHwSqEyeI/aRP7FKSXO7wY0yIo4YR6+wNUE6qPiph9
VO16fzDU+crkBdaorKwGT4hIS1Se/hRlXQaUZOOU8rPB20W41R3BqWYh6oGRfTosxMflGOs0UKbN
87+Stv7Wa04UCj5moIky4+U5UY+GSojXCGAcULPBJno2m8uAV6ohgmhT28SslryGweJl9sWiqwGF
UvfVjYonnMzr655K78FRlnMaw4/jcf1EME1NgyeskR/OJLDt5ADb+vVm5c2WFcOJEZwByobUwSiW
sEnHY6Y/SoXO/ZVcLR2tqXweiWGxAOM4jxEfQDLtePE7Ksbt2O/RqP+ZIc6N5w56nacOQm1AZqIg
emwNBw2iLVKC6dBUH61cP4zu/kywwVi4UUJU71YxUgbcYBRIlizIMCq1kFIuYBSCyq6Fd+tO2t29
vzMAWrElKy0IA9OpSVizDH/FUsYsLdJERMIPnbUHDVh5yWQqWBNolm7tDcy6RVGhL/LuYQDlMfeW
b39pVw0LkjQGTZKqHqj07rmql4qWF3Esk59kBJ9uMw0FSD02IFE1syVjdnmB7sUO0drQhUAkv3Pp
IFS+au+GBnOIcKRtLMnlSx+bPuucLLbBExbw/1BcAoO01hQ8aFy9Mi9/ffqL5kHPXdMRS6mZmJe7
xIwgE9IiGxNKvxiKb+2KRxJmux/uawne45kLsNeaxP1KxdGfyjDu1Ff54GrAvoNWV+Up97QQ0oU8
wDCqRduIk/5sjQ1JO5ZkFLl/x8aKMs8xoJZlmFnChkRp7S+IF5RvkXn69XqpK1IwJzse3RYUcIR2
UreK75GCpDanKK4dQhlL5Vm6dhsCfLpGzO1UAC1MCSOGh28cCHHPPKVO5gmPAUIs3RmUtgBrIT7b
n1PzHtihXHFlWpmcyoPC/Xnklo2raa/2IpGGmPrA/bIo/E/UjcL3RKVCWQ0iY/Ks0ILuc/ilIIGh
9BoJ/jBOqfwc8fne9TzTQ3NO0/EiAGpcVjQd73wJPznL4zjZGhT9UN08Tg8MhU0qb6c3Jw6ufHEz
ckypdWuaL/V+GnfkhHebynEStKe/l9UwnfQUale17bGfIrtHpGHRNceqfKh72VKlB+wf29Ryx2gs
P80H2X5bN8CT+eZAaXp4e8hyq3sx73TK2NWRssMi+J+Ead6jy+GjEDF2GK0qEPfwlTKsisVo7C0Z
PmlSbgX3dk9Snx6XYFtMYDrN0L28g3gICW7bA+mpy0QEQHoAxAphSUtRFBqniyx0heVhCcNzmwX2
s3bibLdGhvddJwgqHMJFSAs1+tPF39t4NnBxj37FmnOVrct/zz8Z/uhCML9g4wIaJN8RaoFXcHKd
KwJBYppBT+YNgRQJsSxnbEya1HmZ7Y9JXqmjL0Tl/GcA68UgPfjh+co82nsPbYzTrQGFecBCLvh+
4BaUSI/aZhZUwzlD9gqk7bmatIBKBpKeiYDN62+FulZ4LP43daVVzQeNnb+N+z/AidDQnQKq/JRN
YYoKRiWN/xVo5+pxeTs9niaT/g7Lu4GHV6nvToL5uj5HMdxJtugFX1cWmI7/TwbgTtfwqp8UaFAb
0Xwrvl2J5I1qERm68pnw3Jmj6zdZXhlWwv8+fMdeemvCNr0CZyiX0V1GX7Lb0iFd7hincpYS2V5g
P599XHGMubiOSlcscfv+NqYcBD4ZmAtHnPUMWESNWaNxXY5/IEZN3jWkdPC0hDAiGFUgpy8jUc8X
puJbW+XgzO0rrc2UNNNC+ovAUhgr9ey95KDgpwB2VFCTEvTNuaPrMVCl2F/rDC8sB2f/qNqTURw5
XPR6tTmX0/P9UaHWl/P7ZqlStUB2T9ymacWQV22g8yKPeZ92kBuxmoalTcIWxvmjZK69urZCqkJw
xr/KdtZMebX9Cbe+ePjfNNRMOlRsiq/sts80anAdzjXRfagDF2s84+nuooHjXxKvM4g/FZ4/doST
Hg9yxF5bnlyATI81MnNuy+XwQQaeBvBXzW5e0/y5/WgszpaINFaFeOAVtEQr36m9s1lJybQOrGis
FuTM/zTcLxcrOqWFeBqKCaDCyzJx/6qj7wn380soILjpZkVAmbI5gYZQ6B5eKpx9tG8HtQv3fRv9
Yf6dQoRf8jQOCS3VLxorYUoxjzgtKTrWIGHabW8iMoTuZ4HA56P9+vleCLnmyFqWPPC1x3Uaf4Of
w5tp8r61Lhr52IlUKPjT6UTJf1iGEASkwZen+NUHze8qz/s1SbRFRx0pHNg2piV9bVrmGnMH1QUE
/jc2uJKnJcjFQsWMdXkmAwPYdz9yJ3cFX22drbS/Qod4APfWyBv4j42Xwt/NQVJi14SQm6WxXXzb
l45DiLdK9QMnfGYz7rbIc1RvyIzdTeFxrBg0sid7+FrFNVGxmIoUYX2pahS1x74PDpc7FidAkqOZ
UiB/aGfOwtPrvM6icnmatZUPLW3UflR5+KUK6iMyg0H79k86idqyP+PZIgJmZetzQL79sZwz3FbU
lMVxDixai05jCyj3eneyn1OTfZNPjph5vis+bPhzKUg/2vGTT8Zljmll9opRd96fuXOwTVxBkmdb
oGg0NDLu0mV3OrxB3P1cVKW3byhFlhNWAznH2zOijoL3aBeQc5zy6Fvqw7N5bjjobYwRc2f+a/dA
epg8AR0u5s0L8uSijvmXK6L+oaUbRISJmNpccbgeAu33HebRNs+iLE5Z7OK13JFnoj/slRQJlzfw
Z4MWN3LOWWNJreBnVnteC1SKxyhKVs5O0gwm9Q4HIZVIcPkEkogKhTjlpNoPGNLztjQwr2l9P+U4
q/zX6waQ0Uv71Ogz3xKrw/OgcNI5BLBoX805bkEg9J7lKmn0D4I9OTICe5LCkz+USkZNBRy+y6sw
OPpYcHvoVRniKUk4flQwpG+YCFrQrHv8f7QdjaTKFp8r61f3XGrUKfFjeTQU8CvCj+hlK2lH+eGQ
SK6iJtZh85a3RUgAx5sWU978mf0GMY03KIHTL35B2kGovMbADiF81IN4OHVKmf9+haxHsh9jvCE3
jjT65tD5iH6OZsfNd6eacAQrXccIyH7rgJ3Lmm3VmHfTa1Cy3UGcBtr7zJQuZyWFtwN5+A+S8Qk9
sGUUrUxuLm92LJJ/VH4Jn6rf6NCXA7qgamD8ptcliKziuNdQ+tNj72UVE7yt295KJDQTOQxfubCo
mHw0i4I1KjQQr2UZyyC7XKRLwcDxJR+zOc8oe7MtwatQUX+2G7Xjn1XqfqR28RU6vhWsrtnK6S1+
fA6bBZPzXjPOxmuz8cQhS/4tBRP7ifPZzy3QMrF5HY0llnum8sLzE10GeUs9JqvrM9g5TNyzTcU5
+tbZxMK+xkbbkB5x6YVpCjt7tlYgeTLVyNwM9zp/4ZlfnN4lWN/9RJIB4cnu72j3CZmhXhQciRA9
8LOhBtl7Zirjs1ddoC8tR6+/XRy7Ff5wYpEyFp2yEbTNLGyduBe60rbfHxINOMvUPL5qtF9+tteZ
ZnUXdmZ6xVnJKX3GpGIbuPqKLuBzWXveaDsusUFmc4pFdt2CxT1D1UJzZX9oxgzIi+WNMVQk+/bW
fAk5CIbzJgCtZV3D/aSO0Uc+NECjgyNTJBeRkwBzFpSaeoFzDSAS/ZP7DVQhkQ2GXFgJbFS1hsPh
diqskVC5lMEWBAOOvsg1Jt1Ciq7qU3sRY8zihFIFUYiSioR1IHT9Z7TWKdFpCQAfwAdwciTHF9lr
6nEx4xDSSlZISxGE9FVIoPXu5wv6ZtTQwbrBanC4LgAkCuR1ursJp+7E1/+r6kK7KHL3geCL3/ND
P9r5scDYbEIX/tG6Dn2A/BPRvEitKphcyIluSzY1KHUgIBWXL1ML7tJbvg28/sIBR4tMRjcLbc3U
Z7htrbSdwVu0zFtf0YLFMTPhpHAoq2kUWCXvleIJ+VZMAPiXaCTb8PcpCa0cAomb/3ldOXXOnXJq
w0D+OaHsf/j6efL0ONeUPwyoikynnxRiKLro07eH/NvOV3z/cBC/z8L10sCFoXCSgQekSQ7Z7t91
hp09FLqBFjbTqiz5tqSjPDRXxJugEQPKHZM3Zar+1hwGrTA+ajHfL3PjGz/oBwS5kkrjmRIFi2yS
FkZQncwfY9u9oT8VHV3KJAg0B92zSRhzK0AMWBFTru9mHyw0m6tPIQLwgvlFvcqDpod1WxDl72kH
p0jOfTejMxgkXs82khdNFA2YBFwDpiu5bnx9+h14m7LUQPR6FyZ1elJ9zWPTPphC+VAwlqeRApE8
wO0sZuzky+OMP0RLoLj9ZhcA/8G9gHsicKMDa+bECZQVpu3V0fzFQOGuJBxNCexZR+ehWb5/sxwN
HN78aZdfNuXcjzf4mujoo/Sk57t1vBfIJqCUniQKjJMicR0639mVsLhUf5FzaQgSLqzGLVey9Zld
4O1huYKDiPl+nLcyMqeIY9x+d7OVB1hHj0UG1WTAWHH1FszFH8VVWiWu5ug6Q1qirqMO5xhl7m2p
IRUArvK+dqC4/UkozEWC7/4cGyXnR1TREeplBXoRZum/XmfvLmLwAJdUJ1GcQ0REpvbkuP4RRdDs
HbAO5R2yn+beGUlNxVJd3pGOL7Yr1Kbe39hvQI3S16pOBPc7wyo3dzWeSgLF6oza9hFDIVsPWeLg
+jNThi0dqtMYFT7YtdK+GQ0vy/nbGUXgQYI6y+Eh5+oDTrkufz1FYh4KIhDUTuLb963B+oOFiqJr
XBQEJXTvkU7pKDDmGwd2x1xbj0nnW7r5rci7PDJMYDlfUcaEWDZzjbPkF9PTROj5ZV81Ry/1Ifas
m87NY6Es2zCiVxB9JPbFsmoDXakY2fc07G7jnpvthdzrqbkODkq1m5MTbR2KwfO+DTmw84D0Hg8M
JDLuNEcuOsmDTIK7nwFVaoCx6IUSTiHtTc38tIva2VBprRrAjbDykYzTB6+oOKpKSeg7XVaL/cab
sqH2PPB8iphTy9uZqVZAg5TB+T9Fr2e4nAeDz8Y38hPOwruD+SnON6I8p/nwfz/msrcQu7D1V0YB
41RtwOYzUL/gmMFf+9WV9upngpjZvqFBRaI7PTmgn3x/Wo5GwklaBxYps2IXHgA/eefHBs06zh6H
e6x6v2HXjEzuOZ0mV4M8W97NClmxJpq63bpyKmeshwZdUQ+LGGrE5BmtOC5ooNMs0POgaghHbMoo
ZmH8lSbQKv4PwQ4l1DBCfLxCViZoHytQZPtqQGJeomEpY/lumCeiaduT+QIN1j99eV7sdFzpL92+
pMVL3tr5cTKM/1QadH8x/jWZHIQJR+qr7/u3Y7hv+PySaoYuJ/75cr3/VlWpO3tanSemWOviUtmU
TMQmqQ76R5vivP44TUBSN88RRf+Zdj9JqJpGFc50lksSUgeLvqwIdScUy5rt1oa60Q1fEJsjAqCf
2YTO2UE/H1tXJZIjGW0+PwLdHitL21epPn92c9OQWC4SOoBcpw7O19Fsccct736iVCuT530HC7Yz
Aj4dMAZbbE7L0tkrjj7OjD7+9MeS7i9e3lAYCsuEe1DAWgFkEp/WKrweTRKoOjnXQB2gNjMonXvS
w3Ui20rXEs0JYeplZHf9PuOTnVQ+XrD9BzMnWtDCeO0nFkG3RHeWt0N3naFEUAf9IychyT3kBiqx
IQwcyBEJvu6rASWEqSYLDf4jGcViPal0pPDFj0mQLERs/U8U4MQ3As3CISgdZb5JawRfOpQ6EPge
rqsnwTvlpBRNlGJcL4vu09vJCBMla7k/cRVGLEQS0b3SvFyS4YiBGwHWbkxhTyhCTV/EfXXqKmyM
BEEiIDjX06RZPfl4OUCK9eOGm8tQPsbZobQH89w+TsRO+J7zhTCdr/FgX/ToMphv1m3pZXM6vzcd
2RxbkfeDz3U76G2uGMX5xk0sMZi/OLJ84SjYpzjH2ru9MlKV4KUlGAFP6tJ66EzBC4HpiUK8egAH
QHSvLkrA2fHPZv3+7jLHOoaKH4Vk62L+hmsR0JdHXv/aYyylb7Cr4kI65cOh8T3wrKUT9+1tdcIO
MKjpu/30+7qJULyr+IdMFbF5MG2m8UVKsVLu+h7YGcQ9GCcJh2lQBw1r8skjt/yS3D+o9e/+kRMz
bsUSNTGbZC2jOeczQqrJpd4GLTYGLRby0kwPyi8Iq5gNuSV5JUzzWZfoGtMsyQLZycMR4puASCdF
9rOZOPNg2/MZnIfuuOYPQkN+tRTUY3Q0Qc6e1estR1DHAAPNnNPXtfutes4z/dmGb/Pwx5j+eMtU
5UEkjUhGFUW3yVCYY1qjQCnGgd7pvkInEPDvOhlu7bo9I2hWZ6v5WZfSZJazPKNfYyk8UzbeA1w0
a+Grap8j22vNVXPgp85pCHsALlz5FlIVrMkeV2piwd+0pZf0c7FRIfVx3gS9/JCjFPJC/7dpueRS
B4bZS5BKYhjoaubbca/+R4Z+biF5JiQORz4RteMIajnx2HkIfU6JnRtKkHWI/Bm6bVztJoDA/OiY
r6C1/ryPv0EKLku+ltS6fXRMTM66olT2ZudOne48zFp6Fdrkpjrs0otRIaJSWOzyE/G7eu9hMuj2
TK5z3nTPUBTXaG1QBETZwHEDIDDr8dPtG8+GxJlYJ3BLoAAgQZuFljD+K0luHXet4m/FvbWKjrtC
bBTNOwKhx5XGomwY8Cz6ev1hLXHeVg88KGUr98NnevLC/rvfNbRECCiO5Os6xIS8UON5y3aXuHEt
hhfZ5XyjTSKo2M0pinuD9xuJC7vegd2HIS0hJ8s8cXYP2FMStsMH0hUnfw+zx4Sw9LofyMTuT+Zo
oPsJirM1DQ0KgXFntdLQcRlo62loX6vhuc1FegPtouBaxx9aii+XWlQZEokAfLfEwnvAHX1q/qLw
bXApoKnmugaRio7GOXdlZa1LZQnKw3kjnPK+Z2hoDDR5rVD2I+ucbO+9w6x+mtoYPn9P0g06y8Ms
VXXGVDrSTGagw1cE/7WltvHUrXGo4vtfeg2vIiUWtISareK96BQpbhFYwIwjV2Rs7KRfAp/RAAhZ
neAJu+6iO1TdlHrtZBEuyDJG78FZi8MFhWtQL8sdwX8glmicg/ETwYVU8Sm1sbpQeoB+klV6gGqo
sZvbT3ZLLsejqiqBbDXwHf17y/6/EnkBfRoFI4HMHP5EoWawkq8Yx4gau+HHQ5nSjlbl5PvaaSTd
H0RWRbAHBf5c5lu//zevPweEYQmiK51FHx5FwRH9dnatwYp6Os7JRP6ztGAfnm5LxBCF1wFxvcw2
dxbaJJjcXGNAhZzmN5ds111YJFt17guzgqG/v0t3ie+69mUr8MdsZtb1ItdVK9dRQo0OUO3tY22g
Zr2VKq03X5srjj0jsD35Pdvu6A04vf1RkpNkCQEhW5xG1xvM6lUtFIvJAQZb5mfiIspENV1sF8rt
GxlIqJXwMAeekE7WmBUMI9mTq8YBJAFDt5Pnd2bodkaWnmIVnR5Tk6bbiGu2EnEOR5SwByhKsAWJ
KexhN4YSkDb5ZqydcmkdWAijlCB1vrkN0Un/rJ8LZ5RBnu+1wDBrL+2y1a/ZCX/6hw3nUSRS5XzG
gJehigPYeElLNprvucvDN6au79sSydTwDC07JD8zVtrjvDZAJRnEexkLOh9IKsci8+vSI6gsMeNB
tHeVX7Z/BmvzsXXTxb8c22oLKyeF3saeCePeePR3pDi5C+OCLslIr1Ew+6TvR5gVCWWBp/z1scbm
mxMR4OOUaieeNhwvnx4Ud3O0sZb1nWokiG0EC26dUqo6uWPDCPqjYGE5AfiHGiidlAWan0mwKf8i
10RdRqHNYbmWz6O2oCdAQ5u6l97cCTYI+T4RJ3KmfGUbNh/Igk7TddAf+7x0MJqgprFxcNPxvmBS
bNp1WXixSr6S8j5FUxfFdMfZTba5RUBF06ID1ORHySKqMBLxazHO0n47gL9WJoGLW4wRiWWuzA3R
IBiWUG9CA/kNAfauqRwf9SuH7AFcmlMALy4z1YfCUhSTrWHv8q8iA3t9a6MXU80Wli4UGrlJ5Rhe
kiReDHBqo4F1DtXJYFwFar1HfFgZLVUv6nz4MVjEwYnkyA0KornrGgk4y5G7pRZDziwwhM2VxQaj
DQGWTVoKu68utz8xEzoYUrZqHmJgtm+Jc3UNurgnjUuFjGOGQlQ/evm9d35uCyKHj+SIgZHkypFf
mLj4ePPGBvIXXyiGP7hn4bCy/145Mm47kYcEvlIxiFfcXijpJgZReOb3Sqn2eJxuyDWnO2y803ya
9nTIvvelZ8pW3SYXg3VcZ6WzqMjp2C89UUYrlVDBUOUxITK7IbWgYKFYqZAWw8DGTk0Jz4yLP7Nz
0wakxiT6cA6+J2gfpPLgUnKq4HMA4R12Edx1uWpsQ7u+5mmmrqEDwdSgI/8izZ9DfEel1YtNf20I
OighvPknQQar6MQrjN2dLfqWO7WN23lzywjBRJMp+p/MdHU+iySkXyJDEGN7TS/NYW4cmmH0h1K3
nVJLBxt6etBeeRagTOFgRhOf3yeaBH4ZA5bl1oaJyNBDiJVl69WFSwuV6dsBErlka8WcqwnWOLQf
j5tEQ0nk66IJykDhPYtYLbnUbmFh9Jnh4SJKd8Jl3Xh4GuitW8nxdmeaR8A/PLhFnYzmHrDS7YcF
BGIEd5XqR5wXxVxiXQ0yfIU26nRBdSMVKu/9cTv7s4ntJ0QV5g8bMGbIC2C1oVDsBd6krOaXEwPR
gwX2zKWrtNgsGeV0p9ywrOfgREnE1hMMxb9pT/IfZXktz0eTg5NVWXbCCQ3jS0OmKVldtmRiHqTr
FSNTLF9htr0YOPf0/2EdCq3OzakuS8xGNNlK6affcBhfg7iNUteodsebusfO146tCDoqAwWwXeFD
dys99QgxcWeEYB2sIq7CTTL/+1jgyvvP454i73LJc3rKsI74/+UL4ea2X9+4UJJ2XRmUTvDF/3jn
veYhYiqeeZUYAk4TqX66xmBE6igGnBzA5DocnGd8KQ59qFXwnimtC+XP2VlOOs0qrCrgs/xyNRWr
R/htRl1yk8+9WluCt0Hg/D+uqyG5JwtpamFzc6gHAvxiJY1cpdQdKGJ1W3+fgepKE3QxYv4ekjpi
pd8XIcV6vy2YgUhNTUGV3zeFAfcU6q29EmAlStejWw84fJu626r5KyXZVUM3KiyF2cJ4bjX6a3zS
tZdZAdUBDGuw+PFJLQF/u6vR9X4diFtHCF1jq+vfb+pKBnK5kY4twIymTbaVuJaQUmPLp11Dn75D
jq88uz9KaacJwEi4/T4jFiztswcgYIH/pAzG3nn+9ywGVCa7DSVKGOF0C79p7xeQrz190tZpf1f5
twxh++9+OREiWtTL4XHHOTRHpS84ymEjn3k8o/vFEjvfJns4/d73CmjI7WZfzBuVFL0t4Kjod0oN
0kWatA6jM00Yzd5ffGXugJKmpwd4lmBW3n2xN6A1JwVGjvly3Xtdk48rC8lCKwGSeN7OcJ6GdCbE
JljpA9wPMpJXI2jM6mcNkyuKWOKoNtOun4qU8nUEHvZYuIsTnLZWSsE4hp6NqGKswEuB5o5MRqep
ZHP9Khp6LWK6G8MxIsGoHBMkivDsLsVoctgiF2ZQtC0YFOiDscsh4Uk42g3DofFWEjUsSGom29oQ
gPEiD8qNgIoXW+u+l65hcKv7FinLfs0uAt71DdNzNlUakLu9ZqULLB5tT7uCngQNt81M3Rk9dPzC
PC0/Rk9h98ENbarRc6+yA2MH3CaijFjzr8WDdJIeHkmh58JumRxNzWGqyv+lhupPEOH8tdAqv3n4
usmqeZgllGbQOZnVmWZkr4mKl+u5dtxuF9FRzSlHKwTJnh442jvH5WLf4iWvPEZe4CzUprZRz3TH
fYxn2QeHbXj0+SapCJ4Puop8kR1NwL6P01qXZ3AUVX+87d5WTdF6Iygpy4mx28Ox3EZEyuD6oOwY
57crbP/9RSIqYAjtB4o/hY0pTmOq6h6yVuzqwvlaPGLCN0OF+3gOfULhae9DChAa/OcmWIpnP0g4
kQCsLsXUniPFOjj5Hm3NAo3myVEDMy61Lm+dWgQPWqVKV54vh5UiCQZOyK9lLxreBGsX49LCl6VT
rFull+gklO0P1rQ5Jd55OSSgAbpWa0KC6pOvlze4wZ3+5FMtTt2apoXFMNUwL/SJ10dpV/n+ggN9
/kisJ09ZXCNmzXZ+ejwG7mXDNM1MwVc24O6qTsvgKnevoGJhjShnwtDC2Mdy5yukgzgrQQqNVk/u
JGHTZIYfGPQuEDDjNYKh1Zkhc5+ZEi11S4Sg0u3G132853fKNFx/O6ic47x1fkhFEY2NmZnjUcPa
/61yqpm65R3I7YChdDIsW9e5Jp83UpKVtrieqBJsNcuopSa653TwJr3CCSIGsaBopAsa3w+hxD0X
Fb6jhlcVOLMH1udLrYxOjX68IuE/FwCoWAMQljACFeV2pDUxVQT3XQjpaNSau358qqpaMyWW3An4
nrTTVHJKkw/+x6CCxvrTAVlWWvl/OEdV2PYjyRaf7v7b3Hr3DPRGBnJNhGSmJWyfsr6Lrf3nivmh
ORkRy4bvQoKzSr42Scvpn99BogCSA5njXgtDtaEZAPND9I+zueiLs0s34sPNzjuCEYFFkwszUwiW
oHW+EPyPJdpcTRGPfRcwhx9pwC2ArocTrZDG7CjIH5I4z+suDvg2Rnpwe4YV0PQ7kNap+Lhky1Uu
IRz6LepuNntDuxC5YjxnxxaMVXPxUfGKJFSGGKMoB6HydJTWPWQP5FcwP3uqTeypsdIwBGy4Yfy1
8dw8fmR+Zdep2bFqyjpF5IbvREOp1yFIHrnvYUC7OSoIsObwPT8DbNMxJVtPAydlCVMQ/vfsc2I0
AROAvZqHYBs1PH0lyJAz4gKzd36QlszeN7ZkgakHedUiEW3IY5PX+VP7oHDXCQrQv9YGS1+RpTwh
vy8sbujDym+JPR/ZNzjLORpWJBTyKmWLqJA170y6ngAA+fdnO+B3zq4pDiqkObU8W2uuyQowBctJ
3LevKUUqPvyZ5sZIfHZMHjowzIqaMU1jHg5rrDX8+uZcVMJ52f5VPTnChKlT35Ajf99huJe0CvRq
bqCvGvtHtN67O/qIUr5iFEkvTVBIwJLzyEZJe+juEuYJeHuaPQp1i8xasOPL2QWoCw8jOUKEieXa
0xKXaowH2NXoLoW2PreVtuVfD/dhAYwpDagLY+IFniTWjuzX3yI4B09yAverXbqVi8uiAdeX608D
Ay/OwQ/gnLhHg25LAuwy2aIcXG2WY3RlFT1ewur+BbLyA3XrdEPQfRcnw8pzHZb+o4UmJPuQheAa
Io8ETMRRZw9RiMi9QL++R3y/X6qex3HuSDPQV4nepcAJaMJVdOrhhT7SJasumFt4AC/J/VQSLFao
c2wpcd51xHadoTjm86W/ZjSPmA76OntRrfV/BmyjhC34PBbgJG2e+4rP5k93ZCLrchWliRBfUbUS
LdKiXVMiWEr1IoMPk+eREgHc/8q3oUldBFDL0OmIbszp3dVUDnbqyjJ9OTqfHYnnciSUkdck1zB+
eNhtGgSgBzN3y+qoW4EJLr0eTb4QS5EqvgAbLr0Iphy85nWH4WrgAFHHHPWPqBM2n+2Eca5/M0e3
NaEcMjqZk60j1xBxoJsvF9FFYYwItdYdPCO9Lg+E/EdZdI/xznTyhfdsx+pO6/ghBJmnLjaQMakC
rxXxFlU71bTEFMMQS4tvaOrvQYEm4v5/aLJEYdWVebRStZ3eG4zZYg49MrJEC1eci/NVhzhREIne
M7x3GTapOeKAM5DKTkQx1oWsYpR0jVbwNO8KisPUXok9DR/YrOCtZaOaM1t0pA6Qaj/OGXDjMjgW
jcbM9DtvJy0A1TbHaMdvx/6eH1druT6fnWN4Y6fXqA3dSDYUKE1eIOM2RjHrwlCtFfL+jFChFkeW
3H6B/AREdS930noRKrnbcVEVWFZ4WtO6J2PLYvEpgyelN9Mpoo0D4po6AZF3sO4dRBvIvr+dsXzK
Q0qD7IcvsGv46GYC6kFLJuwShMWOXMVeXqA2+h/nvEw7TzRG9XJ07tpqMtpHqjY5oEe/LO+L5dko
CedLCb42CGDibJLF/kGlrddS7v64iSiQ7xnBEGBxrMld2dyraEYL5z8xfsxBFXH311XC2X9pxprn
MGK/7El5GLZhER4ABd1wKl+SbY3wEIF7Y7ULBS7TZGOhftf3PEVOr3iyDlzfIviZzUv+WX0V6z66
eW5zAWJcqUDg3eN9klGFufQ37tPvPO3nEZkFlGItI26UsOx9nqbgBTmpMXlkH7G5Kd75K4Bod6dD
EFaSXv3Sf1xqVSYY6gmWSOCsnOQQmoGrm6XxHD7hHdCvio72gea1/1bD4sBosrKwVtxUt5Sl/2uT
GpCWzgzEu0SNsdpAyOQu83Y5LYGOt9NE9q52Psun01I7pSpoB0kIE8Aus+o0rqVdcxHadabk8wIz
4lM57eFj87sCJV0GJjgh1Ssewy3xrbF5wsZwgQypLU5hfb4itDtQQIbHb0sJIoDCxiC7UloLp78A
0Xfc7ZYS0GbPB/k1/DsmHMCDL+hEMPvSXofehTt2Kc8X6OX/dXbfqc2oR14kMH56bk0L8A4WbsT9
HloSMgdhfQDgU30Pw89G73V3p0hKH/rXsEgIB6lPlZzauE18yGeFniSm8Z2tHHBa6GtEeug+MUVv
WRFRll7qLANZJJ7BeLpw/o1cOlvQ1XFyjVLN8FXbyuyt272C18yPGz6w4kkS2tM2GmNKZzr1J/OB
sVq4TORnaezCVx24FMB6YdYxW1ShijS0ZHG3CzPk1o+cTsRSD2oo7Xbb0wTQrEwM8320rt/7m+75
4JQsG0d3tPTxDVP6mUF/mas3ShOklWNxGCUH0WwLUgljaAhIB2EB/tRyFRcZw7aMxgsoQAvs/kp+
m21j25+C8toBBtbmqq/L4YaW7UcD+T+yaaeTCQK2lL/bcqOHUqTRYyPrCAyRXzOfPqUF4mDew+rv
o+Ksumyg3n2G2jS59Ff4naL6anf8AsOU+wBNxH/U5xyddbnRMvoQN2lVCgEdWfEasdhkl35lDu6J
wBDHx2ABzT05r1Wr88apWY/m8s4v6GmOPYnJ1iBbC4+WogwQKz8Yku0anwPiFZGm7iNCHVHONgUp
dIw2++dX3TQYhMr+pc9Ynaczl488s7CLHYHS23jMspJ32YJukeLn8zn87Tnyr0+f3X/JCI+P2GWp
C5SZmETjhlbrUcT1TiAUQOPdEB+gHEnwMu9hjP2ZW2RShk/lHf5Kb/nUtkTBik2TSTB2Q+CDRX7m
IuEGd/PTlia8j2HEK9z92wMPol/SUgn7omPHrw9dALP4DRw8ulFWuHAc5iHpJEHYdk/Hl/6JyKqH
r95+wqoLAaQNv6vHUw0kRZnpO73443vbLEz8hMBM9Bq5BQxd8g01yD4bK3k3RfRf4M7UzR/M3yuj
LOvnLT/4ijXfVR7S0eub6z9ebio7roMjC1ocJMd2VE4jCIUwFBeNwIoPC57MATQEBNo/8bmS093O
WK7ltQsXhF5Z0i5kqIQVg0JNHgxwpW4EXO8exqBbh8D3CuA3tSce/HtknDjwBABm3QnyktELvCCr
IzLY8C2KuGNGF6pg1DStWinCqXHKFpMxw8a5TQc9LhQ/Prbhhrj5FWtUgSBnLKKtFHh1ypAq7Z99
WVJPw/B3wir5ZB5uRtD7k8doCEm75JVuqZvgKH8kIYeftbXSaRnlNfjDnoq5zQXVCDL5DSwgV5PL
I+J1zNRtNIvxRH2C6WfH0GxaKw1MCE01l09hmX+QwiFgA0jGn6brxoDxk5S8/B3/L6fqjQRirGJL
3m97gOt9S4Ek7kR6UIRwPFMBXdTN5Wenh8XyvauHywBp3NNd2K1s11qxVy8fo/teqAIM5/qXuXQJ
GAbdZdZ0b2Q+dKc08LpbGbDY/eCeDglDNKJWfRLxToJhBUJHUqWFlSS4ala/t5CNjJM2btTqGCSP
Af6wtwcbRfS9Xh19oiRc1teC9Pp3cegxaExsJS7hjqOI2Y1tDnN5Z6G/+S898F5vwqDz4e77z3Yp
sO0Tq9Gg31f499RQ3W0X/xDrp/wC/Yh370gb1dYu1uu7c61bkkw8Dif4+uOYitXk0Wbq618jZCXp
msyNXDr2FRF9AGBGSZTQ3dKMUjNB/aTcaX73Wn/eDz9woEAQ6xBtwapMWmoPc2mYqoo42anRFNkz
JbhTDPy5xN0Hn8MEcye3EqhfYayncZggMdHZm45BQo1Bs9U5c6T3fQXxNAbYlrSLCd3hZHLrI1iM
zTXCsP7nIrGL5wq5enpbJb3U/mlIGrQ7fG7bnZDMdNFLPhy4u2ncWjmTYKDIzK/SDXCF3BYUiIaV
1SwdjR7P7lNtw5pGc0WPRteiYM3M86Y/4nC/d2xVUdFuDcCt9BrxehQ5Nlo0pNg6CCaIF9et/5jJ
uCptV/5G56cXrY9/q1jAJrKqfmuPhGjWo/wLnhIB3TCtZj9+FQIhHZRVi7Gmw0FqP6bCiB7Ip5xI
2zPSIVSVqYPnhWehEgt6r7jxjCyjcLiUz1UIrh4ftF6pi163BCxRp3joAOXA4+iU4FpFgwSOuszE
ajUvq4o8EnYUyt4sDs9OhPJYEq9UmCz/6mR/uSZOaZ65IH9r4Pjdf5fBPesPvkXElZ4QUzALLh+U
91g1zkD/MZEsRZhzT5/KCf7Qo2tYBT/Kg7vbFh0gf7wq6cpgb+KAd44KowRoqOun6dxyktF3ObHD
1TgGWqy8FGK6tC3Utql5qVU+WRNmR7LQGIKK0Nglu58vz5uj40WGQkq3v9j2Uh73o3lC6ddVTLpr
06UlggJmrYXFhyKPrYKBFqkPwoU2WH7czmzFcNu4nMmTP5z89D40k5CvwGvdVQ9bla9gJfItVoj5
svChywv0XmJS3ZvzQkdLHN1npSz0jJYucrRvU2F6rAv+yvWXtsAysUfbGrgvuSiXPQrsIh9J0gGQ
dFgEnapO/BmNLML2ydd+uwIIQuMyK+S5ncMYrnaNfK8fYHwmwqMFwJOYOz5WrPvhhaKNGrW5bdBH
7b/fb5J8EurFl6YzJ6DCvdLeRz83m/bxjG0ynh0s9YLeJPFX+UBK6CBZcy0Sf3raB5AFIkybq0FY
9Gh2IF3F2XExMkzxuAsIbjmh4mBdgT8XHPFY9aPhRKU3LQFLO+JMt1s0aYWMPaAm0nLrcYT0+lgK
CVsgYDLY5enMGev/LyvPUIGUOCyFlFFR4V1dGkhy1ze7yG+39Ys9YGGKiNQjGi+aCczZDznh45dw
hZwi+Y5WCko+4tdBWSpJ8lYXcKL1JPNXZ2e2nc1mhNYgEpzqGF7xU5jx3LePXMZUxCZbup1i/htD
T/kbzS1Y8D+u3ZHsOAFK7S0hLyR8g77lRH/Tk4gBs1Pi+JNkbhRcY48ZKJfcGn7KV2XqQXCFynYi
JEjORYUo27hCTXtrcvIJ0Q2WP5hIj7FovN3Lx9JYjQGqEa/VmkW21mtQN4Ek05Uc+wTbUc9AQRrE
gRiuJw1iExVi4SP5gOPfcO4nxoHlpAUo7mRL257lTuTDQX8ivVzkf9w8pRjFfOPXsftl3cL3MEGu
a9phCplAyaV05D2ygk/ZOtC0FbgP8CzGYE6SFK/gP5qllXHqTnHGBq7ntrDibwmTkngl0QtUY9ZW
md+N1KhWEM52FRVd1xsJLrw/mqPLPiRtwkxoTBDPMmcnOhfhDpYbjj06xlsvR4bCPKJzEV9/5wjl
MXdd/0zRIpUFxFGRvhccMy6FTt/ce0/6cWF5XYrb2qd8mjnLqg28weOzL0D6nhkUfMRwW55xK0MV
cBzlNHKk4eto5869fBqaAG7qvIRt308Dr2aLWkV8F+8yhrB7J1Iflm+0p6I2w9Ip1/er5d/ggoml
fUv6Wi0zgvBRuX665p2FXCn0Dl9eGvhyFfxPldlpM3IKG2YGWB/sw+mSXx1leKQ1pWu81cDwnytK
TsDEjTJctq6w8Yx5SLjTkGsPoFzKMjI5hgdWJkcjvC3EA++8DGb1m8+z7EBVh1LIsq1ACIcdv5ZL
Q9UBzxck2GDe7eTEoYsYOd4ohtHHJTuV+fVbcyMM06sZcXMU2st3YjXp0/2I9Ieb8b61rhTa5ZkM
iHGWVsydwc9YFUIzvF+6HzYib36iQiAfduOD8Jl+KR6GvQ8g2wCmdtA45w8PNGzBb4xqLH3wgVv4
g1QfppPQK1THt+0AzVr4h6ePZFh7SH9HAr/Qr71ke/k3jNLf+SSaY3CzcCoY+hyWkv8RIU8LYjpo
kRhObPlR3uiX0hv/JV+VpRpEbQLj1wKg/rvZaJkgK3ezNoCrm6CxdRT6TugYezBjnh5e3d4jpzwr
EXU1bReGNKZ/3yS16a7JdLftqJEtyWdoQpqSx6pNYF63z4hyAmVFhfERWIjPbVJ+DazBU/PUBCzh
I0xzmCFvBwkFFbPgAdIHK0Q4PaXwQesuoEi1DWsS9LSslwN0o0kRcI+bolLInHfoJYONzoTTiL1v
iB6AndWJuXfE/s5oi2UpF1BE32gwyCSZUjZNBsvGBQ3ixcl0hRNa2JwdM1lF6EYgcl2I1KipmlZQ
P8EsRWjF5HPqcu92wixgjWiajCTe+zfFs4TAKSA37MVHhK2Q0f7p95jM0Ii9pd4+jQgEVEhR73DB
mTOS2/K1Kl9wdeoN5m95TYAA3voAkLLODKdd52mMVdlw535MiPzttjOeQja4bA6xdSlHvGMOqQLY
FCBBJCDyrTMDIP+akllKiKnLgIOmngpib4ONS6lWOtL9rnjXHuHXuM374IubM3836kJ0R9vRbEic
aHUt5WRBEETDyTXdx0AMmJueQ4TyyxsJl4bmxNBmx4CtQKPXXxQ/iwVWaL0ygYgOQFECzJbL0Fnv
dleduvGLj5dpoNmppCgC+sO3DadTzPmtFIx95IrOW6N957NjFK31NirJ06qcxhZ5JMYpA77n5/te
JsHiD7LZ6uSD4261Ji8yxqzSd7+VMRV21ArncIpTpw0zlMF/kxq/iRXcMwMq9VAOoKCWNb8QwdOO
3nVhF+OR/c/HVmEKNs8cEWEm2I9rGSRGtJY+9bqtoyakArhs2SpOn6T71rVYDtCc68wuXh1Yn9y4
7EtNDwDQl3WVx7j+BEyANxIuOF9XuVOuGKRCPdTqJdg4JimWK6isg6DzZ/faisRgNY3xRB1FcjwO
wxRi4CYgUaYLdnUxGPqMUHSH1oVjqOER6lok7R7rjOEg8kG8DDHdgB3z7BXIzTH8HOsh13a44sY2
zEfAM3lMLcHR9YDHL7hPGcjWEN0/WM7It9XWTKw3r2Tz3xRxumwKODLrddIyzB00Mojx/1vDZnDy
kv3bFYAuUp3ftlFgjK9oegbxBfv8hhEBn6AxXx/6TNLWYud6Gi6L3KDJOL8F6rSuxyg6L5KCbIkA
dK6uaKp+Dr16ZvcqLBr+NVITAwYypi/u1Tvn73dt1wv1sgDmjnioUdfeohCj7l0WZanXb4Z/qwAl
efIQ6fnYvdO1gQ1dVSMe33UiTWflA6X43veg/jdI/Ekikk+0vBHCST8eJvt47R2p6BH4c44XEvdd
FrOgT9TC86lJrrpgCMKJci5AP8wIoXIfx0oBktbbXAMd3fmDwCxLUyNqI1GmDQkf5AoFvyJbOGQo
WpVNzcC4J6Nvl9gWpOpFxCOKM7MjqHgrjc74XzzXmkc1bOog4QfKYh2XQUGcjlcN0IXN/lMcZCxG
01CcQ9lip+Pz1ESks5+h2PA2V48ydxPl0eiThm/TGR5cu4i5BSWevFiHRL1Kxuq3L3Xwa36D8ZM2
w4QygqP7TRlYHn6uJIuJQlqqKXadKrNjjWZ3WObwU0lfwvWmduljwfQPNP49cCjQGsReR25FXeF1
bN34FjQMGqqqJ8YOzBorD8CRXDfVbSycrn9RR7LvMpJf+SVkLZlzKDekKI2DoC0iYHwbs1J3Bv+Z
gk6Hu7g1j625VKnaR5h/svqpe0D/ziqtOmTr15nHMLMElPwLZwwyCfPwQzNcP1hBWP2C1xzbhx0u
abhaLaFPhQeAGhGCN9nlOUqN9ofR/G16X9LmVgK09bS0PD/FSI38iKLuWTRsiZPlj2KbEK9bX6iM
pyEFMHf0kw5aUQeZ35pcPJc8B5MkmpSV2pbpRYkRgQEKxZE6CKWp+nA2mTrNQvGKYVGjy1FTqkqA
N5aoikhWSimX/q9TAu+j7wVVS4LsXBrM1GTW9FWZLvjlqksQPWOuEkTYLJbJWaiBEBSKfqNa9220
L/M9iZWm4EgbBmxt4Xi4bHTQX5BIdiOY+zs9Hqa36WTOmNtMI/qTyCPgnz061pNWCMv9PooaYy5f
aupMz0l9qiy8uHW0kYNweIiZ/q8Wa0fAOEmTIdD0KIKD6FE/Dkcn/3V9K1+/QVCSOKS2UFUwJYrK
Mow23TZQ1O1jlE5x5D5cqSD0MHePik9p3tqm7TfkIC20CsIXP5hmSBMU/7J9XoNNwfCysknBphFD
EVSgCxcDdecSj2Y3I2kuYoALHglWJO/egjkrFtWgvrShxx8ed+OMF+GJ4bsbZtD/XKhUTRVxHAY3
ZHNTl5Vqy7d96mLXyQggoGtdrZRnsH10FXHA1ai1tpo5DI5QCCczpkTF55eRLetewzRenn44SCn4
dfMQOFBCXS2ka2/hxy7l3aYQ3R2I/8czOmtds+wY8bSvEVRFsM5a3QLeJMsM4/xSFm5OQRaWHSnG
3ZuOKHTLATA8o72c3NpQRCHke2n7Z3HjQc2btNGfKcM2ujCxZzo6B1F7cGAy8NwNy5YKG2pWO7YW
zYuUB7dUysE2utEb6Q3Fhd85RzpZeIJW3LbktSrKNUtokX0XJwunQol5G8OXszV3bkn0FwGZxci6
fTNSoUf+Yii6ofcuK5iQL8DqLltLlLY3ORakpiqrRRH9z8BAIkPxg1Q+vQtG4Y6dnT9XqWWI0+GB
OEZ2TIls8GE696mwhhKtfn4DvMF4M1Tqt/Oo16xEWEmKkmnCUD6WtYmVRKknlTY5JALpdj98JHVj
X1NcXzaK10nYjH40c4EFngfz3qBpfVKcAnryYbqpFBN2imN1K+Wsj/IITf/7shma1nHVG5gwaOje
v41cVYgY8NOSvyvjShE8teKEWcdoPEClNhe9vuzIDsaiXzQ5LVXIFA51YCQbvXtb+SUnHWBUPilr
R6yZKF56yCORuRxKT716lsu4Sxy2t3W+mJGLIfRp9U3bLo7blgQalhLR+PLh0k/9OVaqJoB8z7Tf
UPpXvD9vRTeYyBUEaHSzILBSFuVJ2BKUNFnXukrxJsw3aG15AeHmmnEw7FkeSO15F2Obl02iodQF
4Gh44dra/Y3f7EsaPojP9F1ZI7nRO+wc+VHvLKvoW4SdzDFk4Lpnds9ECBikgp2DrBv+IC4f0VR+
FlF/pjee0t3M7nXDNk8KrxwgIfolGFvoHtFqeJb4fRAJVHoDnJKWDFukHF4jRzzkkW1GIm/DIqC2
5pGxXMxG/PsDIZ9jhkGvF9etFIYocpwVsR+bl0t6giEed1P/nnMusS9Jw3zYa9kPgQmRtsNurIXp
AWaFmKJIzK1CQZFKPBgAAhUVAQ3mHOEDjAnvr9OqvngmkJOzpSrfSc0hH71k6+aNoKAXhmPF5eAj
5b++Uftx4LTtWmNvAOlTAzXbSzCdfo4ttny0yGj3G8y6rdznD+k6me7frB/db+iHxrvxxY3GMWum
O93XxnbsBz7s7tIQFA9g9ZgbfR1f64Bhw5VRqGaewrQ/YriYF8j7xSGwvI7AroR296niTt2UIpfU
fZ/gNGzCWLwn1sCvwuLLiV4AML5iyp16Mh0s/rU+LjDX5bqp8min0a3EUjO1upxz7DkOpqQ5bFvS
i4mDDHC7/KXjSfpvoiND+BUx81eBup6QC+Hn9USUAccH7hDf+Dz5hc9Z7XKHVqVFDxVjqYcSJ7/H
KCBEzCrK0vcqZAPetdLTm+hDL/w14yh6AErtbCBDichXxPekBzky/4wok0i2oqs0dDkoCXmqJS1x
EDBo7xgnkLno2eo8XKLl1gctPfZI0pwamcgcHHhraNO8+/3hVznMqB0ADXzmb8h1yO/ob6L4+7mD
xCcm2sxJ58jtOd7KOHb78+0CYuWHbh5WN+TkR+jJBUhx34sM3QwOEes8KAHHb4nJgrxgSWoVd57F
I/FWLpaKiAQcJSNBaxIAU2ExyJaKMp1ZeV+puMbWgslbIwK2oJNJDyePR2SBDAXV+HoCzYcK0Xnd
b6IMBBdybVDQsIUFpWUDG1O01i7PnhWJbCKSxv90+un1gJKw4jTTtIQYyr3rZMmlKsnl9+8Swya+
NWjmvIm7FOqmz69ta73t5Cl183vdtlsO8R38GLgo6IJNp8yDHQiaxESL9z0ahnpzOQD9VUkxih91
80KaOuTg8lDeE72nynoCNkM8TPqXTAl8h1L+fxkwhyjzDaPgWcEgSuPTmpWzIMCuP8M0wBbR9Y9n
uxoaNguyTC8g3MdvxhK53s2RW+nlUF8NiCDTXCSakIt4CUXd3UwLVJWxvwwPkpgCSZomkVl2gUkH
AQ+sBH9OgSEK5+RQVAu3gz6AEJPnACS6eWu2aLFWTEuSSAO1bUWa9CdeIkTErdD38F9V12DdMHdw
DK5rPHOJZPqPkG+069sUj9r3ZkJU2oY6FwaW9csqHUGdFHNZBPypNxDfcimGSRa685XL8Eo4SvDm
zAEb6h8xngB6cnOt6Z3i2Xcf2m/O7BldiyPnFncD/MlRmxcwlM3MW+MaCdaxTB+T8JvOW3kc3M/Y
AQ6KV5j+xRr1bE2C0U10iI9XPYLXnQLmMG/2K3DXhQBrIT4znCCPe/T35SYzkkkw/DR0eyW5Ox99
GFzXsJoNvw5ZSE+vZirOkcE14TZZ+tuGkwo36eoOPQtQC/8gIWEhg5/A2W2eIpfSpC7sbARTslge
C3yGy3U00z/pKXTvRxYN/JgsEqY7omHbmg4FgZQF0b9WmE4qU25GqaPfMNJI9Pb9VCEWBAsag9hT
rAKpqfmyHO6zIQOXTSGJ4iPgwgWwKE1WIa2tc7aTdXo1gDPjc2mvzytHSSczTcyBZz/4AZmKdgI0
fJYgp05sclZ6cAr+BHlOK2BkXMf8ZnTEjL02FK2VeDTEifgmENhF/rCnRHI3hMl+wF74xZXA6tBd
L/lqrikXDR2377DvdJvHBPnAvUFYkaVJatjoA0s8U0z8IUuJmvrU4vfjUz08tR5WGAc01KJHdXpF
1/7/rKc2Kxo3ekHlUNsSMqBBmHGHF7Balmtjk/tT39Q6n2rNCUiBtt2TsJu6CsGnGLwuJzFzNmfn
7aVGsTm+TPbdbNhz5fQsZbI1QY25GbDlehEezdAMW8YrZvZwc3UezEDcqyLW7MD+BiqYiz1UKiwt
43GxOfQlT9dQ2PxEc7Ppo7m4vwPIgLnrkdiGxGh7oUWGOkIJ7l6wYKClJijTbitPossAZnJWm7YF
q+3uC7M+jvvWxQqmPFR8Cphte9FlxSVqoBqCHz5wR18arjuXNH099X3beVioZZXXkNi2MVSECp2g
EohLJyS8POwhmOnQ4PDxH2R3g1dyBT4kU+cUAnh3/pQW1PgEJpUk+3Vktv4gtLW8cN6hEZfAOlcQ
dc8K5hqIZkgb5KpAXsJpuY427gQcPTQkczmgJ/9CbVbAIU1lKME5vraCEG5g1O1e1233hFOvYeQA
Suqsom4HbLFCmksodHNuihWX08uo6SKQUn1OpPuNWvgqPOgXY2XTXjl2cbN5X+pwsKC+Vg9Mow23
DWEgBDBX2F6RML6Pq9sIEpbVT8u9/MsASDzOXy0kxuOpH4MzmkJCIgKzCb9zUn59c9gR/xTv7UDS
20lfx4EwnALUTglrNIIAhUzfSyCJI7pqpgKbtaTWA/Wa5hmbT916aDA2aOAEwryvHWgv+NO4ef7y
q66ngkrSKuwcTNpUUdfRAREzljeut14Ur7KQAOlw2ZKyMXZijon4kWPYxBvcColiMq8ylzLorPF+
JzDHdVzAzQG4mNsJhUzqg7vymlu7hFj+H/kolkI39B1wbnAS/Q9WoOSiQdBt6ap70yEXaokcBUgi
JSCI/NecN9wc1Thax5wB5WbelyaUnvnjALBUWYaHodyzEC/8uaSR8h/R6Ndko5wjhV7Q/wOTEALR
HmrAkk3Czm0jtqZTC8CA/3fCwMtrfwNt9bFEFkAdJ1hsQDo0tDSsoRSXQGLZuE0b1AxjuJOSxQrq
1TDtbbCS1+mFn5TIJpjfC/KacdCxC6IuxbCJd7ZodHAK0T8vlfL4X6Y/fDxRPCCMBXU8fN+oXX7h
jbEMCr0wwiRz83k01zxQ09nX/+b2C4vx17Rg6G1D4ByIPhI9wvE5kgXgcsAdYFEoJukLeMWcmGwe
ijmT3E7ksZcnZ31bFkl2v4gkdpk1jESztFlWBARczyvxyxu+qLBwc/O7D+gdSFyaLn9rc1T2vElf
ngrR418nwuc5nCZFwdiaFzbCg1o5SD7ZCuUmCB8Cusjv/mOeVFpoRAd6sPbcgHfgeemHO6rpme7N
M6Y24vtJdNwjKVUvoOUNfeSAUYz9FBdCrGeNnIrW0TjwmrCalM5Ii8kgJi1RmZvdZcAysvxWcZcf
H3owMSJhURhkde8Fve9ke6fGWOzsL+z3CyPd/uK7O1k6rvHr/zdIw4So2x0DF4UefyUQpfGc5IXF
ftUjnGSx3/uXcpAGyqOYDjWA7WMpz9KRNqXbQME5x1cryALTKUSZ/wEZf7QTbokhkHBAEpOsV73G
8AdjKAqsWLm/fZLEuFKY2ws2BzU1zFT9vwjTmpX/FTpEfTxN3evDTk2OzVlWOz92ln4PCQ5vEvUB
bJ//vU+LoTiXKaJQKhB/iCyrZJije+VgotvjOjL0Y6bSaaEEBfoQraVwCGAaMCBVmODaRS9Lr6gF
oXPCduQltnhnEu7otyOeZN/lzn25ZGgzYjsc43X4MwcQwOtW9m2ST/gFLssTBZUxSxB9F3TusT4e
JO2KFoD7KJVpPff7Nvft03ssa7m+692bqYIxb9TKiLLUOqSI/EDmbDH0OnUQWHcpi3rLzG/Vz2Cf
YO9IfQ30fufiEq9U+xQGKnopbJtbLRGzKCRlw3fka+FjhoXXOmCL+J5ZMcgnBTpRp2qpw893oK2h
fLCIDB5MlojnlR1fzSpvkhQY6kiH38Sz/awTCCqheuxB/liqb8DQQckfzgqgXd/nj+5vub7Y7ur4
LJ7jwS0/5q92zX9EFTdEi+Hn7W5MPYQT6vqABY3H4Ga0JS9zVJg8UrbF0EZZzwwfRvjRf4K5pzog
1ajawf9uakZbZTeQArSYNaoqnK/DDOC4LUTWS1hGLMEHU7eN4OaKAfz9CMnJbemgpgKLP58MAXM6
4tji5uO2hvcC0pMWPYAMBNxomKJFy1U8ntt4ZcGwDvVW24PxfpFOc0vQwatMOLJ0jN/dLBjBkij3
NDLAHm/XgwCGuAzl7+0UuA62dwKsusvhXvOvpH96XAel4UkobjZi2HakmMT44Li90pTUvOzfnw63
cGBorC4fCx68pKnIfc4defflOfplcqepHAoI0nDoLOomi+tNzWyHA+a+pEo5FccbrHoFBLHA+UP4
/kcieH6klPS7Pkx+iF1yo0aFbYfoJPTvGdyMC0FhOeBATRyFzcjrlplAFi+4iQA1KeE0IuiSDRkm
STM+PL00ugpu3iX7W54HjJod648zg4R3GmzZRCAYpOhe4j4yJXNt+ooTWfEHJds1vKvu1zxRNIX1
cPwZeXLZC5IhrespyDmoIodfsYKqYzpfGGL1gkH20f0SJaPI2IZerYzHT9CXJQlZWmhFluzNm/tL
AWQMhEG7eriE9M/J9qiE8tVwHN5vL/oFXH1s9rfwvwBXNc6fzE6bvX3+Kof24+n90sscV68E4UGY
1ir/0LK6dekHRv0PD29dquG1mk41Cm5IzjRQdEjyWHh48BORticSm4QZ/WX0jqQj3TcY/zEZL5rC
xmno4VqDEpdqyRReA/Bm3174jZcCZfdxmDk57EO1U4FKHtu6dR9TB34VoEDwqRWeDzAeRT4kiSae
ijDxFwwayOUxt6xWaG5Wj00joB681ZYl3nQxlzR/KkfIPWUKGD6IwU//k4V23myal09Pg2ovBmH7
91f+VNB37lR6n/5Q5DwCqXQC+6do+LULTz5CrxjkTr1zeFx5dbeASj/+a4i8vcQSdvU1bJ7omhsN
OF6Z/x+O/ybO0OLA+fFAlvhko9oyQFyWCDLFuDDT5NXpY9fC9OAUPB46wmTkFzlzoIpw4rcXW8pt
0yoPOBlUydLXezV4cuYthINMiOinEeSBDdZK9/UNwA0xSkc10nQNCtZ/CuuEG0HXgp9ScPWwMhYL
AYU1M+VMQvZxcalE9Jy9nZKOLzYs+Sae04iVQPSV/jDUuSvq1cNMY/M0/oEdj+jI58zXWk6WqikB
Mui8Tem3kPlUbRf6lo6QblKasWSQfLsBvPp5m5sFmlutyK/t8XF8OQVTbHpokqGgEe/yXoQSSl45
qIGCasXW2gTPx1BX0KYt3lNUiQEXoURlrdZwp+q0mlEbDnn4mMOxqni1QwnJrbo4lJ9CxfXpZRyC
4UPZ0OMuIiIDh1L0skkDF+36h9NuFkAA35Bb/nmGzyghOWDL6r9ZjgQTyxY3pY8HSszKSnBR9BJT
KCk4b3zfh8xOPvuQ6TBAmxJ5i8p3CBrgZ4Jbgkc9hshx9HOaIOzzXzgONOPS6Xs3mD2qKnxNYDmM
ckzeoAbcVMkAI4pRxJ3WuffTve4uOCiIQ04OqzZS2QuTwbTRMGJTSP2qoo6YBUAT5jXqD56exAaH
mIgdcOhTXgvI6Zne+uSsOT8A+PhiqMciMUluRHgxvSy7K16+0fch6kVVa7URmg9AtYMaK1hPja/J
KwK5hauy/iX6TGjdW5wJax0+//VM45u4XgXz6pnWCVI+eVjg3oD1lW2aVOnykb8v9rQ5xSK1FcFK
LtzANWm9TDPLyejTUWwfePPRpT7YiENccASmmtU4A8oOxNM+EC8H2lYrqHEqUoE58+mhzYsE4tfY
eMC0xYZ4yHrLZJoNAggIv/gIp2CMsUWnUazRp7V1POAzbQufQSvzNRFp4noN3Cj5Rp1mr8rM8jsg
2mXho/GirY+14lc4RY9Y1PdLrxH05P7KyvNiKj+w3Z9RuGOynLordiwY0HVV4Ai3dMadulMscesm
K4AOAdjy5+ZLlcK82EF5FfUlI/crFb3jjkcQgtalQgnjdhe5cAWRXEpQa4Mvrc3vktxy6KsX0B7W
Yc0+0Xb9Cy9jjDeyzQ0PQTPzWsWmeU7xBgLOTVC34lRpeJMj9b9MB3A39CF4W6pyUPqUtjTNMemL
98Teqdj9TlaI4ZXRUjHb+Ac9zHe4ohUPngelex6TFGtEz8T/fCk0rlqaroIVS9UBi3k50GBSyGqV
6VI9N5BzaPWHDWfVmJQwcBXnXgVNotJShtqu4v5p1iCCa+PkLk/xxiDJgU+qq6/ISBxY5z51PGHZ
iI+9JhM0k1o5Qr+1Xvsah9AKIQJya0nrM7BT5CTr6QNZipCiTlcuV9xiig8vwLDabBefsPbIFSey
Hc/TkrTySj1eUADuqFR2rVIBd+t7YO4EzhWEg/K0RjOevMSGI7wwXd5Mw+x1gpai1qnSinZ47v+6
h+bkTAX2Z1wP5bRU+1YqFAza4T36zCvH10lMZDEI6tenaJ2BsoYvx9NRggvtnktfJLp3/R0YZoYF
WiD2/lQ6uIczJjrirJCrszdl8vF2BhDjeEooj+N4jBawztOZZZCw4v5riyTSloWsYygOJ0Js73qO
I7zGEVee2cSYlkM7h0ngdKAuwXJyJanp5F7GYDeqztUjLkUz0kA+WV3OoT4GnPNmTEurmlxkIZdl
BrB7R7S0mTl5Qts+ONkY1eOGbADm3C0SYixWgJ48k+A5/ZS8E86YbQ7Wk4vpCi7Sv3XKAaq5wY5y
BHV4qsUvC/3QPoF3SOnXRwQlj7bRooqqKxaWoFX472ZUJa2xfhdwbrKM1AqiF8TPnTSH1fYObgvK
Jws2zXfE048UKY9ysYh2NYGkTMahBznHRcCl3SBO05HlPkcr1hfGgiFYMZTp0U+HpQFWM/EH9qc/
yBYoUa+jK71bNfopEe3H8uwEjpqZTOueKwjlOJQDaI3pR1mD/URhvZOvmOWolMIIZXlthVt0XclK
CDwpycAHTFj3LQlMyNqdssmXTxSaBvJ3tBilGigbSqcA3xQJPSJB2MPe7ducJsy7vZuKTSJ/Hdau
gGxIOMv+IUL3gKgh04p8IfFap5POFFmUzSPMPmKwh3wu+hICmT8ZT/bVLxVJWJbh9y5ypYnQ0jbX
czcZUrYahK8tNrK0h49RPhc/GSAa6wzihGKDskVPdLeP8y/YVVapjfPKO82dhfBlUerZIafnpNee
/4fcuwqqBOZAQR1LK+39o6lchUABgeDU6grMuVu0wCoPj9MHlCTLmrxGXyyIfgA5RJxbP7/mX5Kh
3jta0Ci/LOr5RoH/UkAq0H0egc8fHLrCDNz06wZMnxoOuNCV1911IxPe93a9ua0zKx+gC123A/Ui
rvJBIP/xPaNUHnhOQktcRggPFeeVVyAsl45JLM8cVxsNKbH7VtuENjkoklr1uw/Eu2Gh274jmfpF
bNxsqBgpBAbbDjeGhwDPPK03PrmahDIjlxUTH9Ogvco+SdyYomkhiBfwWycPBtbaOz0tpzALVboy
Y9RBDbJdEjXW7jvSFu0O3nteiaO1sujnUoL9LFXtlYdZ9Es3MS0ieTr6AGuf3HewSk62nYo/qzIS
HIgeCa47rdrFA3IR385I72jGbOlNUB9o+drDnAKDxE16+3GMhknbP4z5GSrFIvvaYCFikF5+Vkqq
mZGs+yJ0TyBzC2rdg+oQjM1ZtU9JUePSDdFUqeIGXXPYdMrL4lEoYg3Y5685vGJVlzW2NxSra1jP
i/Bel7ybg3yBSuLp7oUmLft1gjMjT1b5jiZTJ+vV14WIqt1lSavp7yaSCwe2OAm+ZIPjM5elexwL
P/IOXtEp/s74vjjzKSg26/WAv9NKOT/hB46SYQY6Ly+JNogWyZWJwu2PMK+Kc+syymVRDNqz0k9j
FvPRrpUuBfqHqc4bbShIhqM6j2HE01U2Me3XlVl30dJvQ+zw3TZLJodX7T5Ghxv6INuKeFYaoUvD
H5rnE+74gFqQeM7NggSQVVvTxKHYPNtP6nKirB8+TPMV6HrzM14kvfnqF2Tt6RZHQm0o5zUgyowI
0cAHw7zi+c/6Xr2d3XIJ5dGBaEaaRdcYeF56s3TTNEl8xdxfEkX02dJ6LxWM8+2/Gpj5BfiniIRT
RL/a0egonMP/J6+dVPd9/a0JJ5MbEbimcIhh9Zw5s7PbfxCFeUsfpPhqOTvTGdhcDVnRTq7DQY6c
wMt0C0+PBTPKmsW0hvjJoXiyZ35jHpO4FoLo/zMflrRMOH4qegNvDJlIjiQMbx8uKkwEZ98181DG
U7Bf9JXHp152Hm8hyrDGX1uJpubB0VvH54codM0Y20IwdJ/Oa7K7HIcCRWkcrqZJjRsCEWZ5RT2r
CzzeggofTDj8pXxgeta7sRM/+cZ5PkHxujA6QGBZgwuGKIpesULXKdlj/gpgEgR2s97h5xEO9q5T
k26vcLakE/A5k6XRSP1giL0Jh2Vj/pbGGbg86PBXfA8/8futxwCrUcF1xJa2Klyrw/g8h5Z7hTSn
9+J1uGq3c2qZvshKfaEd46YV83apgDnCTqEO/E8XH0dVFTkG127QLgwoIdMHRi9fcIsaV7zaKhL0
7UttoKhfCdS1S/k0L0kfTgI02s24g7Vvb6eAbzadxq4yOumk5U3cak8xIvqFtSn3lt25VrFaFue3
OlfOyJm1nEy8QZ9Jx6Hzr6a1Obq4h1l6zfk41esBPLZZCfMzuBm/lqpCRs2RaQxUeC+5InNYVDKI
6RDvY9B/UEule1byB0Yco9/48ywvzkeP6+3/OvsxTZVPEolGSKHHRj+PnfqeKSxrZ5fStYtoXBvE
IyeJXjo/2X7z+bW0Ou6vMYnUqE8Pi6834tybzx0d0dIw7aMQfQlMSKtXFpifh+Zee6EfKlkl8LHC
QtQM6RD/OtpJCmfDLpdCngdqdUecNKDtJO55dMAQoOiu9In7pEhK3d15kyZSUwPwI/qXEHMK14ri
gNnrhHSdHH7FZczJKO3UsrVMCbl+SA1FmGu3k46rNoanvw+gjMNlQt4rrKcM/Gnny+pFJPCbByJS
/1tafS0glQIN+hJkbZPR5gLpy5POlLwoFfz1a26aMUrYwfpjKKPSLsj/jeJjoMJmR4kv+tgo3uQ9
jpGn0q0bCGTPLL10sNhrl4vweFnvW6NyGwR6dZ/caYNWjZIT4LYSZ2OsqoOyEFmsz3sepDBBJyMT
acMV+Y7nRoU4LDgvAbSrwBz0VW9oiqjAiz3+jU/mDuY3aNpp58/s/xVlq0fDF4xs44rpNYuWyhF5
vepVbNjSq8co3sYWeRT9vNB6gq9CCsfBxo3FxsbhPv61HHbwGimvfuSp3Xwk2waBomhuFl4QQRWq
VORQArHTP6Vldr8OpvffIOVNvlmFY31/67yaF7ZCkC86oK8+J5omhHeYGq/gKNYRQ5VFCeKt+agt
9QfU/NQwSa0bl7tbmJULzq/5t2QWpdNrFiSsBNwgHPa16E26BWAO9n3KxFGyThIIROxgDbNRy8K0
l0a/3bTTi7mc/itRNnFcx2vZMfAY2kphEhkZmjJ7XGVOTWf/7B5O6wNETrnvC/mXHmlc+fumET79
vuBkmpkT3qhRm2Uev1C8cktYJXEnbQfGh65zwY+K8X4rnMXnZxLH6S3tILo7y7dt5Uia0kHBnFLn
aWHc4jzACFCTmzymLM+GmfLTZEi5+vYUX3uwBi0rXueFKxhxJNHYJQ2QqH5wFt16phyUdkVTWklo
OdMDlYY6D0Z86ZuP0GU80/I1y0cr6I5cOr+uQIot4D/8ZuE2A79vA5noQe4MsgPdO5p5wDTOMjd7
D9IVtz+UwwiWXjoy79LjsergSjQ+UFYBiDxiyKPXPoAxyFWdVHNnO2CSs1CqTDW9MoUZ9R/b4co4
ozzizxN+8b4ddExT/CdihvKUud5pffYgEsEanpHRk+CA/qUzFs+J+Dfk4JtzsS897dv8//LZGPHJ
bCVgpNoyHk+oPAQNIfsfXI5t3YBcG2g4BGPPszE7ntg2q8PaX45PFQMAAEMzPAsAkKzYmcc+Sv8m
+hCkRRJplrnBbIGZbJTegy3bJVqDmYLlTJrJFhyQzOJGxOzWMV0kx/Mkvc+fIBxHjAwabFySL9K2
j31hfYQ1M/CJab2ek03FnpDGDeDWezYZGdB01qoonySjrnmGmr/SUBEgI5opUUNESsgNbARjpZWT
pLBbxsyKiN2FCaJ+G/5p2yT7NHk7c9LcERuTST8B4SAyMw/O+7fZKt65s+LMsQ1CiVWdCgL7DRoN
QZ5LUVWUaCYhFJtIvNwHT5SFghrv4pZqdjv84WBsx3Oy2PIAyFQYDKoKGUoqc9++wVuTnDyINDJT
Q2hBxaq0muWPGrpxWylvT//SR6ayhHC5YpdR457x3o62zr/uqla53uM3AXWkf2tbQYUz6w3L3OTf
l74OFGw4l8bY2TYO2WdNPst1eY8mScdtMjNXmMEnSEcevl/pkHUlNRVLDmRW897w2PkJKcL4K7gZ
+M4l9/tIPLl2pefZwMB374KaeQAwauOJNUKHOjU6KykIcY62LfAox4EeK1+rnwegmEfPZdGy+ASd
+e6NboWI6OCTZUbWatRp9UKaPjTyldzUKy2ik1dsOAj6tSg8Mv5Qpwe/ffsEY3uT0+6Dw1ILeysk
yeupTDKkwQ6N+VGKDSy23iQwiNBUWMvLp/sI8/miBP29Lb8Nk1+V1pyvrjoCiByq8XrQ1T9qbB+a
LofSCWXb+47/DkCflSD2k7c5AzqPFp4S3T99f6dbhMqI+Lnf/U9zeFmH+xf3DmopE3yZkgiHeP9d
KWKFN5EaGlMIX0VXvjxozRItUCwfgMzR82H7k/3DGE77NTbdPzFpF//JACmIu8gdqZJDM980xKJM
w4uFu1XBeWOqjSrR8nwfEstt0fmdMHwb7cQ14yfYoNjLbf+9CN8ilP71E1wEOFlZA79H/J7La0cN
5eKy3b3vhal7h5A3+VGXfq2PKdQJmu6/jCfa9ei7msT6JR/ufTxLXwEQSdV4YDR95Z6m3DHqGyAa
KpwSy9CWHosBZifAKAyBvCjUFBtR43+nY5M8H/dLin521dNicL2xY+wXh0SILY3k713emVd3wUjP
3z25eYOHzkxgl6dHj/4oQkp/4OjL8HwDQq4CH2TdbiRkRhU7NwG8w1RuYp11Pie8P6vbDsrjU83+
mLJV2rD6qPlH+TWLX6rNpBp6XGkG8LSMUBz98QNnph82xmNv6gn3ovpDSy8TN2mLtf4hie29iFfn
7GHuKrRQZKuorwCz1XEMHFPe0xlUpt0TpCUF+I/mkuxlOQez/CJJ00gYqQRAxE4h+WyDZl19wvfX
uNKKE5Fps+H0eW+6snJiHB6KQyKVDytR2rSMcyKfrNlJ22VjItxl3XwXjwVoa25CU920Ku66J7pe
IapnrlMhHdheJtRJw/+Q/Vw8gT4ftzau/b8NwIdrnxbApbrxjBFV5Q7p8PV/zYJeXgi6vyj1QocW
DgTvk3KPJpBUmcbF6LjCu4UrH40C9AmYi8ZBNp/Op6WNE8ulN1Pc1DamfSswxPXGmQax3EnYL5yn
TnxgY9BIqUBzuLfFvBHeE6wrbK/3ri2yl4mwrVF1Z+jAe5SKvae9E/+nFqf6bwri9YRpVLwHjciT
g9bugDvGPUA9KdG4y3gc5cCIapmBkD9LENzhxbTx0G+RxGaMmxABj38leGxz7fdwrYqO2jZ0oSyF
v2dkB1iet64Sjuh8FqKAblHhUfo3Hb5Y3CcrHH+jYDuCPYEkGKM81mTypwR1hF48EAEBY0X1fF3y
39boOdp1l6Wwo7kam9vMqgxCC0QfuA2AtaJC//ZCxkCGJdDwgRJYMbJF9ZvJjkmao7TrrNUtDOix
hoqDA3r4ClE2mjT168nxCucWvJ9oUv7F1+aJsFOnOTY/YFjANnVqmEs5MhCR/1rplsXntDQJj62g
3W43pXLtCySz9gBcZafiVXpdoCGqq3ekvrP+aGosWAlaqWWQAGf7uhDHlwiFwvig+vjSG4ETzcRD
yW+qpvcFcST8i2fkpuT8c64dnyhrx84qormZk+UnIA5Kkhde7m8Xk/L1fbt3YzryrRtoSTxhUNrw
6ULvgSZvwNrmv6WzwPmQKycT2JfsdHUiJaZIeG5m7XfQSVmxxYoRH/IbtaSNSf739+cTWDAoVp/T
BrUnwjV41Cor9/Foc71pOgSDeWF96rmd39SNf7fZS/Z2Qjd8mPFTxM8hU383wO88SM/k6EPdu4eQ
0UM4J2DQzTiDollG8kDqSkgExWlmhnauZGgjjN42LOBBtSc/wxqBio53OjqEs/C0I1OkyCxaNa0b
c+l+tCN6Dh/GiEtYFFALHha2d1rtaeggEFYqdMSzztXe1tGn87XnZTzzCyPHV2CrAhonbaDUesgi
KpLdGzYxK43JMYROipepSAQl2hJ/RRwzq7LWIjar1QjkTZ+bKVNl7elm3OSGG2ZJ/xmVmHMLBKfC
cqgMGBgod5Oz9Eukk2hjpr8YTYh0kBu1u7lPnjZSxQpf3jg19lQT93VR8kPH6hF7M/AAZ/oT6+xX
npTlG+iV3n651qqbJMf/4HxTBzz2F+j7ICeNHZ7h+BcYsvGEBOSJEv/PIDFa/9SNiJln0u+mFQtn
+Qu7eM9CUmChhL8B5F6dM1NVyvEKa8m5BqOYXrRGDSMG0R5hw3BSo77Q3xh1HrhEa9kKXLtiuuXG
3uFKFzZsvinwbY4NcpGz0T3nFr3V3RHz9UqjZjBXlrwa67C24cs9xEwxFq62qA6PlSTNDk29FODw
O8/c9LagjooHjQ/p6BKG3+d9VBPPSJiOFthFjnj8EzQSWTaJh/kF//aMHfLbJSPFPsuJWBVQGqN/
LD6X1pvEtR2OgC0RYVfX7l82Qt60jJTBRBCrP8NtsbVSkUN1Oadg+jM3UE9Yy7rCdNX7xwslIgcr
b1WIiacoPy9RGwHnbPkzlDf8h4f4EiIH2skhQBXe50E1v8W5O8969T9eDcr2vCFfXl2cHzedx1wW
YY7sDeUZLXBIHzK+7gFzwNX6WjVMzf7XdL+aEft/JyNFsb4rX8K21PdjIZqu4l84BirIPr3RLSqy
ROLDecdTw+4ENkdxbepjYd6w0GbtEW7RhjDTvLJPUos0EOngWA9zxjLKmOum6kqjxukR1udVpjf3
hO6EQjxarUbqH7QCRvIWiCYk0d3rYWNRaErtzORMOGkcqcEmyjDfctCcgQUAnSb1v9SybnnDrgh+
0hNqWfk2rk+1ZPGCfxu6Z7899bl5tCHIP1KOrQ5HcG4q4bFw7eGgohk0Ew3D4/FgDycGUYYzVIw5
1DyzmPx9Rf620f/lQJ8gjI+h/7ici2ob1b+XgtD3lR+xSAprXh97OY0cUPkJ0kvJxALYE1mEfBJN
m3Bsg3KsUCri+Kv3UjIEh48xepvFJZRVAjmfm2pYYrTYkOcPe4I/eNbjyltsDsrWNzOPis21vUyN
AwSrTFCq1VVpnCrgAwmiAotzt5A1I1esbujI5nUw1cZ6290VQF75gp1P+bo0rHV7nPV/IikS9XRR
LpOiN3Eq5yqA5TydNwd7n08OzbEgw+7NspcgwZo2VkkoQFgvWHP6Ow7MmYzeb09uhHMKzODPZHqL
tma+n7i7IjCh3GWwSafvHrWJAL/X7KUfFVip5dgnpX6wOkc+SKDzAFDiPnJHkNUiEIUus2OThNxD
T29l5RhrCUR2VYA9iWz+IX3pffVJ59pZ1mX/yXt3DiURtCzxrxKKIOFg/c2KY/ZeVDI+kmaIdFTu
no0F84n5wxLqCUSMNYR2dlzoYUAjLkChg+ZnwHDVYr1S51aMEXpkmPYiXOJNEWYtYmelXijPtNov
g0RyGqluYjAGrJYwN6TAC0tE9H4ZKHM7mlmuh387s5rsKywwYANN4WVn6WSdvXSRDKFoS1IEoXLa
4za8TAIAy1LiXOYb5Ex8xT5d3nDnx2GL79LNKizT2dOk6NxTngQypZbOrrqSCa1HG9wOmn+GqFe3
h7+wSmdOhfADp4WzUdouY2CCSpMJIDbG/NTknskxRQkTUGFbbO5lKQC/5ZH6jiA+8fQ4mRLONevs
NoTkucfFnnhhOxHiLlmPMyyIVjIuEk6+JJSBVjMpcybP3L2IoEAV2j5mgn18AAFJ4qjnjCOcoIiV
JpsBX1rOLUa/N4Fj3q9It9YUe844/C0xyCcnK39fr4UKek/PLmSkX/ebltgTfEhmLGNA+F99IA2c
tA2PdkWDOlVrDVXarqXGa8l/SlOTJmQfzFFgo+5Q4yuNr0urGzpo7lyOqEhzV4ifRynEA6SX0N2A
xnTAB4Fn91q+Da9Egy7twkjBBMYjLdvGbHrhfxe9z0FW+bbXN3CkT9omiNDgoY5QfMnpnXVZEFQc
FjwEuYcSKj6s0OLFNHWZ0RfvU4Ppdj+50baaKXog9Cx0HlknsFXmCSAlwfw5RyTqH/qOKE1KHh5W
8Q+vO0uBlF9QPqmy3ZUlBrwMa6ijCAjif4v3v2Rpdmf2KczemiGsAdKi/EPHL43468O3ZV4k3yyj
gr2Fo4Cq5rMsesrfrJEZDa552+LsyRnzTyIzeO9QneIWlYd2FqPSkRCo1D2Iykm8+9nWPfFgsoiD
478o4cWXOspgj1W58ot6Wobzh53LnjP3eAVehiIh1wowYHd4UJhEzYigTWG6AqEnOU3SUbkHaSpN
3cUF5jkLfga2e+JCcHJAnEy/X+2ugvm7gxnyf7sakulVjqkEwuyVpdmweHEuQfcboTbw/Hya5B48
KhKk9THETzHb3yZOZmFxSKF80+ZCBEKA+kWo7paX/EAK/BVk0T+uyy6T6EFj9UoFlIPrdJxNO2V/
XElckzVXe/heLUigk7GrYm0zkpgnLSbPN6dTth4kN4xNwe3mLC2b57kGX6lTEEbH4k7Bc78ODiu5
XA5jDfRr6kvOZbVsM+e/A4T05VOzI0AvtwdFL7GnazsdYw7TsMFCEz+X1ezKnCqQNnPFcCs3430w
J7DXXrRnK+qp/p0ENQhNo82uILFhQIcG/b9Km1kN9xA/+Srau+vWU62UjobNTGiAiVroFMrk8SAr
z24nnc3yyIOJPPvt4HXMQC4IqhSWY7NzyF889hmjXa8yJiGeyfUo4mx1Fwars4dCDBHc1GESRlNx
6touB0GpjBmbmOtZ1wxOmLGIDifaNJ5EbtJbrpAyCtuEWUmIaOZLFyW5oXXyVcV5942qeNbG4bSm
FP3Qm/iQf8S+4+y+nEFTM+eVaydgcqgJukQv6dcXj0GVNuQFViILeyNmx2J1/eVG5TYzZiiYqfex
3i/oT5OgL/Vnk3lf2x+KWegAuRym92T88vcv2hZhUQ8homcP+3yhvoIOBHWofxFQcDbahqMCULoJ
qCkeo5v/MzCros2UwTRPSwh0Z5T9rzdvcDYWAx2K339xwjVilyoQqrb2HmPX04C2YCS7AKttoVXl
jJ3zcoSavhLlrkDTQjRr01wz1fcE/bSVFPUsKOKvjN/GppEnI9CmtgL4o5WkE9uFnpLMASGyyROy
jdlk/d+onTVja1kwcwLIvhP6G7jQ8b2wYQI88vskYeWtAWYL35SpIESkyjl9DPTpnKzTxQFYFuS1
3ZxESG2a1PaPNlKQKCf2NeRFZPO+/EQaQjPCUTQCmDQwbDz08IGP6wMQf/pthzh2nc9ZFcZDgF4P
3n+DKQWdWqBZkb6uIR3lEYIKFmxSJC+DU42Yf1tUSw6+XAy5bbMAD/FAmMoyp7BbalyMYyy4HFsu
u2snD6TFTk0CjL3u6T/6SFbfns+kt1U23xA0kf7vrJRYruApWa0y1xAvbN5yZQT9ELZ/J8gST0tf
X7XYwtUwtWThNqunWKaS0gz1UiSTz5lhYvujV+uekW1NGrt3hekn/7U2K0joAKemRTYQSH2CfEs9
wr1v07oFKdXy+y6BYIjcZFRv0XyKeovMubH+nVQHN+BDJsrh4zzZZ2j6b9Eh2hi0J/JZFg0NlfEi
COy7wz40sIIWqzF58TzDAQmHT43mJMeTLHqW+Vm9b/TaMmRq985KpaOdsWCbVeJ4iFMwMw+PaHYu
1utU7qZARHOJNITCaB8SrbMT2/Bw2HIgOMyphjW5SQiKvQrMwevHJsTlQ1qgkwTziD02Gcxy66Kj
uBjScIbCpvuPAof3uwqsPEePLXEAoEQZBAey77S66M0SwY5qd3ybH8WBHKeV4Z2MwHeIvjAAnLQY
fSBV+t1detDejLbFSssaP5zh6jBRK+0j3tlIlOHBj5int21BMw/9ORJHivvbB58vkTkXSRD94lRS
HVzj8/Em7fdRzL7FXgV0fPUlf6KYoHBnQekKvTwOgOSLUU/t2f6QQHeMHTgvNX78Z+Qfbqy3qiH+
7hOPVc/Jl0VcgywTiG9fyOK0WU4ARXojGbv0MllQViweD8hCM+nHNQqdH0FbKehgUlJItwkfVpKB
Q9IYAlEyWNDUoQQ9x72/tJNAX1KFpPW0Y0uSZIeRJZFme3pANB00sHq6DzNXiAZJWkezEpcpnRRS
58toSRFwWRkhxCC0mhRNzpIItfq1GnTqP8u9qQaaVNqDI703Plf96+2khFjvWE9wtWH4gjZ60F4D
k4bCtgGqWHHsgRMC1jfebcYXFYsmtfaSLuRrZ2nb2yxBOvR/LXD8pdzp5mNm7yeu8Yf+qO+bQKmH
lPxdaoZKuce5Md1ELqTgKqqHJkKH8d8rV7vU26StGB2/4O0aPfTcjpLagkB8GTzz/oRCUvCbD/KB
ih1ZuI4eo5+c9cVZfL8/QTcYbueq60rjmpIctUm9CMhxOHoyb0u3JsvKkwth/PhMVIyX4gXwkFZq
F4q31v1gq+A68KTYFq8kE1FUNumguNZ0n7S6n1tGd3PLGqZCVl3+cvY4yML6P7uTOUGTFUJgThyj
W4jyPAr2D41WszmdZVEN5FVWuaOgTQ8mvg7C8jfG+dozU4yc7kkp61FuuR+1/M7AH+iSYBhSqIqt
/sQP6H68vooPoKFGn+TJfcUBl3DalFIO8aPxXiiPY/MDRGe6caeK3vjHRioaWEvG3uRG6YOSyp9v
9bzrzA/Uatnz8coaJdtTL4U2cWbH8osN2BojkUSrpvYFqXn98mOPXEuC5S0q4L6FJ/BD/SYURh4W
RRu7et7HxBctUEF+DWqRamWQl8d1TexRS9AmINvFn3VYsxBfzZ36bGEvZJbdyB0SJOhHbTWNk5s6
JDalHWOnAgkCwkcVr58sy+yT5v0HykAehJH+sT0OajyXjK8FPl4+9/WEKqIGtzxOtb1IUMOo32+0
3kGF/5VFrBGUh0SWI56xYFPV2Z+sqVzI+AQmPhWONyjQ9ushHA5hTkjIkQ6grYfK2qgLJJ8JJd1f
wHJrm86be1ha4AGIx33Rt18X6kI5YbavAJ7fyYKxGLyh4L1B31FnEqFNsUjp8uxlJqohOb69kK+z
kqN/P9IzTXo+eJT/b4MwuAwNWbYoRBvcm3POeCLKd08XFSnF2ikuIbMDUdvCXT/Nc7AKfkGBcUNA
OjtL5h0/qcNIOtIxI7vlWciR6e67Tn53YR270Vgl+FkrQQHz+Hi/88YjsjFHx8NMiOXa2wPtmsuG
vvso7cJUp8KCEr5D33mzbN4gbgehK6SlTe/xlnAEssiVPO+SrFKjb4MUDvW0UxJK4n5hSileQEE8
FGzOh/dsJH4NCc+cJN6FCkEVMlJF8kcnPYd8AtiZbIJEaz7849nGM7NnUMajiJ2ZDsg7Xp/SbZoX
A+gThDT5yd3rWQmuGKh4rms1j3MJhmBdrXmknTZC6+xvOiaosfciRYSLoW7oAWzaDEq07x6GQl4Y
H0VRasfa1KClHR5WYTNIRDJGgm5phvwa9XqgM6zhesNkvKLvw73zhTH7PRa+IcJKVU8kPFXlgUGz
HKEXjkovX4uVAbwB+wX2Ko9o9P5K/Oqu0IeK8WhwpKqXCq8LWPfC0jBkkoWXEqKnkHjj+PqAoyyo
E/BMl99K6Ty6YOaS8/AFAt5GObZZ4MChd34wN/7a0D6oXABhlXQX2sm+vJOyYEUK9vkfSgMgtDPS
CbG96t6VBbq+fyD7DXniUrtxLyg914o/k5rPbYfLIjcqqiVVMA+YK+djF9RClwIr1is4B8NHhS1Y
oY9K1ofQWTCaFnnqmqDFBw4Nb/7Ak+AAAMsm4s3Xf/QX9KyrhwodsgSidufWr5qlDboqwZ8IDvaE
utXKvVDkEiXtAguLOrxL2ZxOWQ5SpP9R15kbKrLAnxR5iK5rW492YM4yr4ZqEkRi/7K3/GHb/K4L
Aaatx8AU+GbUYlY5yz0St7iwahDFKKD33BWuKX9OsgQy/ZPH6+tqIYAnNAu1NEgoA4JoX+eAOIRv
Syl4IyL2BsbZRhujxqQpqe4Ruge4AgJHAyD6Ak+MJ2f78GYq/ZyF/AhNw9Z9MNP69Pj/RaRtLRxg
NDbflsGHdWGtQKG/rh9y8cyxAufCCk9qBkMT69PGJIpR7tUzpF4XjvPgFl/Ne83yVKXuurj8oTD/
qd9490AXDYjd2I+Gn+IfACH/d0XS9zsMFrpkYz4pLvJBOyhJJ0xjTH9HHgUWvUlf/y2WW0aD0eI7
kDqCt6l8YNoaFedqT9Oe7sglybNjjeeDo9ER4M6RPwHP/oouICtKc9snFd3TDUYbpZuMuRX2RZKE
U0tGxVUvX9wPv5fdG2dmIq2qBrXLPiTxxy9CqnLztm0blmp7ijTwll+OKt7zDDZVFTOYPeyKJYnD
XK0OMkzD9QK1V5sYrFRInetM62rdjETRwHmQ1wVt07sxnCfrJtns4rkmatKKt8Rt9HTLKJUK0w/n
btimH0jyGLx98vgPQDLRW5KaOtTsIHmvBqb8pJDLcrhmbeHr/BqOxq1UTP6alGoBGrpcOJX8ZytF
Pw/Cgs9Vk0o/oWC+/qxtDY0jYnlOCnfDjFQYNkI9USoiV3+JGHxhxPJIxx6nhsg5rJ/nOa8vjX/g
kV5fN3BQmW5u4NCfLCVIvIeZddOBzo2n99te6uZESkXMbHw5dopi+sBh02F/FwAcmuHnb1dNGAL0
uovMNAdqkBVMDAZtcF5ANbKqTH0z55zU9OgvFnI6cb4phksEECALSDELZMKDn9/CxHo3AD5s9AGs
2WXmAXPyGDTPDGHIAVnPM7s+AFktibVcqV5o+E75DSTbUITFYHd/luDIWdof056iohlyMSzurPQZ
jUiOcSydrxfpim0bNF9glYF5riSqyUg74xoekUJw0vmHvK0gI9N//mwQ5MyDKlQRlOey2yJcbcZm
z1HenDoHkaQNhSNB+2dsSxNUxTYcVthdYBonb26kj0R45Q/+U6IwFykRxe3TlXBcR6oGkSXKJWk3
5ccxu1uWs1wd5u8w2tIB/e1nHURIL4pnrt6G5nl7YnyFpNzUktoAyGEHr5zo7AodKgDLQ/6kor70
pzD6YtJJVxe6RkYLWlmNHcKkBw3bwlvhCJarp9+mJWgdECC8YOrFdig2eDNtLp019mDwSZHfxLSO
4kAw1RzunF93NMktBhthFyx51CikIgVsuvwRYhvkwrq7g9WwuFYy0wNhF9wJ5s88N1wScZQ5DASd
x9BejUZqxyeRspxT6obBTTNlJNdKsuIHArGtbjjfFm1mLIH9t+GwLLa5cutPrHvGorQpBNHGdoka
ziL6GlUbggj28xb0JK7dSG337OZDIHX99o6d7KtUsEM349jL6yjRehZic1PEbISKC0TB9UGj7hIP
yOWu40bQVDnPzVVSzYPuBE+p0RIbhGiT3HDf8NUMPX99K6uHV8g99HU1Pm4ehFiA1mgsBMAF7two
nc83VaPqDJ8Kubagdwsng8SWi/K2oJIQwH+ReYtSJF8J7FOyNuHs5IG4bzykTT3tOWt9Cw3pjmDa
kUqETw60Sto3tqMW6lSeV9nu7Selj8QiOuX2P5sLmWw0zcS5zBl+70CWH1JrOYnDYXV2EUGFXB/1
ztsxUDrsg77mB/E+0JCQOLWGzncBUIDtja9AZP1OtL/ZE7GfRNUOwzBpq9AorvVidDcIC3Xo1CRm
65NxGUYOmxHWXRBc0PnlwtdYRWTLpqmess9GjSOJKLhuYDbe4uLFYjDifej/0zbol17Qw4jhfJry
ifuM379bOk1sI8M9nJEHbwCbWcMxn84rX3wXoCVtOKbwl7crzWHc/g0ylQiCMhtyr3sGkdx7qwVg
MLt/lFuxSh6u8ETOJiuWZmlj8JaB+xFIrGdGjp/75tIUZJRr/RKkFBwd+mSgEVYN9jwKAH6UEcXE
mZc08PjqdrKiBkjHMT+9wO9Tkh96n5gYCwk9y1nEia8A5TJY8OgznWbcEpChg2o+aQPtAXcgQMDS
wSPfKncvkYHaQiFJoyw6n+ma1nN3ZIudhjDt+yr3Dxl/TTwEwQE3r0igoelNyr3uSQDM8HgUDbjA
CXAs06AiNa1V2Bnq+IAsI4Kxk8siV8/QPkrxCax0dohFIbQf/Z5F1RzgIxLCD2HH8WCBVwVh3G9X
o1/ThGu4iqOTgKVTktjaof8DOSiNT7Sw/xu54ZRpIeYqhHggKvv8aN9R9aR4h5uEFJqrmipscWi1
U9iTjJPpMoJMpKMB2PU1TtxZqeBleNP929zPo9HLFl+Yti/LONXarWaAewXvvoSiL3I5eGzUci+5
WDiLt0TNYGybxpo7JimFG5l9O1jiUXVyv3VmooDlUpO3G2TVDZ/0rnqMluRAv3Bmes+gd0jCkHqK
gGIvOwPTh4XVNIbqFng5c6zDU713vtmdnggsJ0s+3J+JR6Je7F+bp1W0gqdiiyS6vLDp44N27ETS
ai4Dah3wQ4SMTEQzkosqc0xUJfI1k2UCKobiSAHn69JaxeDxRjZSgDhepCXynQEWvS4JUM0IEg1l
VyE8X8KTiZenJOmDK5vihwst543AfP6j1Rd7WijEurYXYj1RsMUVx6775wFDU71va/2HzVYex8MX
oND41zMp2pTqKwTCfDq1BKx4VjQaQm73yZk3M9HVNFkGLJGL0l/c1xoL1l0HcA1vkbYOgLTum2Rl
u5cqa47XDfPu3pdzWWFEkgeAVXZ03/4KL1AkPgUrDcueXnIkuQvatTCZzXupnmue6MYlBk30glI/
OVqP0uhgLEp6IIqVQ5et/UvXO/mqV3Yz0lcnc9vRY88BtSTRSEXZ6RjhDg79EeTxewfbIhgn+lca
4nBAfDfWzxQW0xUrmhEHDUESYLsIceLYh26B+5C7VEToY3cy+fBmF0ov7mXvBRWPNIEm706Izs6w
zb2oTs6P4esPLdRpKyerIWqzwn6TRrK/t5cI3PAtLvUFq4oCmf9uQzsNbxFhqn0WuMAMSRUiMSlJ
uq3yh3kD5U6pzf/hQ7nShZsgn5qGZ4grS/D92KEP6jjltevZTV/418rCgmRYpqWmT8bKE+EdDnIP
EonaidnroPKjBdAtTwojL2pMGjfsfLhBdxjEg7iiqTEhaEMPwp7rJy2eenIRTOR1Ig2mwNnYd6aS
A92Th3Vgnx1hDmYhjwSBJ7Zb2F/ujjS8eE8vr8+TSb6UCyLNAY8Tp9miTvfheDYtzBApGwxPCFFA
Bd27vwfUCF6fU7rQXkI0173VcopGybwzy+wpZsXZLkzJam+kOZ2hFwdu+yYFMU2Uhq1TsAJIaVpo
6S9JNjzegvP7ad3qV2wAbRIr7sILgWS5AFFDIQu9MY6kkXJwpVNM6gxuWRRM9EKQ9XobWjVQc3ZH
aYsQgHUoqKI+CCgihmRqdckq95ZJ16rXFKL3JBnFGewTlM11fBR+9oNDXi6ICj2tNo6b5+0BeRgk
Q1Us0/nj9DQGLgwZFuU4k1x22sdazdtQQfCwrlAY1wfenYm4sRVKJ35ozYWI8pTOzgEOvLkOUYph
8aRrT+A6N/icLRkzfRBumIIng8uybP6c13d/qRChq5n2U1IuxTwyVnstF67CyAkzES0DYSyhlogs
4VaW30Tt4s6LfIs4yPSYSoYShJ71wiTgRoVf+FUHbndEfG0EMaQozF4zQAPpkBMJog514HfBPSWO
mEt2kEsl58SJqfx5TfWHhhP/jNghS5IJ+Xbw/XYvh5uSrVjluDPuHZ70UxC81S0xyKQkg95dpj+9
Q5Re+SSNI0yTlW+JgjctlNpISZdyy9PfDn8WtEwQfgg4tpw8AE4IrrSpx6tri2baG6EnDWVVKnDM
m+pI0lYl9zKnL0gxsW6xMIQpq5dwAVQalynLN+3cJeb3HeknHo0RqaU8vwGyteV48khaGvR7MCg0
ayjsGGfUDYXV2Zn5vIdzTERMG+5uOgxXqZVGVFamH7sa7DfhLs+0DxjvBS88TevbaZMT59kc22eo
ZmNeHxbxgRMEns4i6EUamQjFC2mkKUKPF/nUTt27MT4ivj0W1vhambh9kXwgdnXFmcx9X7n6Wdz6
0k2F1R/ZdzV+xOfij8By3Nx2aBgyULr+h0o2r6xpWijok72Hwwz5RqLsJxlAYY+okkWWltbFS3lB
kWUPkCmHwDIshsSkcFDHkEhLiPf3U7Wl+nZCQUVmeANTQSGK0uLbGvbdshzkMRjhAggQerzlRf/m
5lgxH1dR6CFlLEXigTHYsVlLFvi5XjhgLRQ8ECJkYtasGU1kQ9M2wHZD4K6fWlD/Dm8Gs1RxxSS9
Vy+KFzzWGNz1BcdHZbdGOm3+9dRkvRKSmNwFLf1S/zJeHKcJckd1JuglwEDzQDdZHCsu26MA5cme
2kpE26qLlsTmmYXFwEN0MVG+zhhDD3cdsbGjx/O/iqZHUCkMA+iV98s4wNK36jLE3QKfLlS/tRK1
WsIf1tvLBsaCVViognwZKoVGd07SbgaOkgjLNd86u5jUb459Y6EQx9EjMR7b1H79N5EQDtzB9pEr
ejFC0HmiepFRan02lzjvTOI4o8qKMlrJHMDV2jaeXeJIQrMXylUnyzBm1jHgMc0tqEZ/TKgbbSdr
jN9HDDQBSdg0CUQtfYr0Sh5twBNSYCIBCK/b8nkda1O/+lPA3PFi20CU4HNPthoymvFqMSm24RtN
PM4k32MBAahyOY2gKHcFLWT//OcwKkIG7Q8VwLkwMExAnn1Ws+4GfIuugR96nUBQdqx0q+O0cYtN
FtI2QdS225FxvKdDN/p6j5tf3hC9uDiHJ98nNozLN/QAd3xEIyrYK10xGZf1MFvLdMQ2LqlebkgZ
7eePMcH7zKiAIfqqX89wf9KTgRXDYLHjZ0VWl5gqUPl1gBCoqebia2SerC+6NzfP1MPLG+ZbgfTE
lHE8y5CkkUxIalVowBUq+xdBwG8RqDJZCrKVkcXor1ZRcAmMM7JTuUScdGK+OfmrAaopsAHnDT/4
3EU05y9ibHVWv/6GJb9tyEmarSwfP4fYmDv3kmi2w0wn37f2IUp/RG+NAVy/KnxQzH7RLYXiBY0E
466ZGldbX7Z2MRqaC2kIAFzqcQENIcoMErsWErTBZ4g19Mx3FmE8fgX0/cWKFaKkSLVsushiOT33
/a5MlS+2waQvPneWn4OBcrxomCsqvjGs+H0iPbsO8mjMvVySgb8I1R8YsVTsAHplSRVsi41P4+l2
qOgLRvqfGKemQRc5GGtoik4MOd4rNbj/S5A9QpQX5/LP13ycVs6xSPhBA0PFGnLi4KEusSRvcgrl
c+4DaJCDdWi3ayUJxv4XXAJCwgKfTf4OrZ9OaCqSDaAYWm3NAYlFNKP39yXSAboJKTjMzKNCy7Y5
v+NU2yxUYobqeddKHMSYr4me86jyV2g1nez3IvmaiMpGVmDOKq0Yf4OEg7X/l9CjXHfXOXHei+O5
USjzVFoeXrZycZYjQej0xx3uJjRlBdQMBxUvGhFqdS2x4ITC7c1b3Jo9z6NRN7hFa/rQHEZz5XrE
WmBN8vh1VFwXWNW6EwwvwLgkikzzTVY5Tu3yseaCG56FBdsvzuN/e0XwbXXSIytbwpkbuUkW19VF
aIAc3CVh1pGRk+75UkFBwjNaYdGU+/DUtI+n2d767qJ6j2tqX4qitcJNbyHrAqG2Maf+/ivyVN6W
gNX7wgewhb/KwtR9QEVWOx+6wzJcN0mFHIwHICifqpDVgCnCEGciDvTZM+w1bImcjjXGdtjZ+gSt
e+Ck20wA+ENd3bjfjsx+7gPDMOoKDafq0d7JL0dfBNMtoDGK2z6VPM9N1dyuuadnOLobdwLU0vY/
1Ac+hvoc9KzOh6+mQv/FW66rmRHLgqfvPL+MihtJqlsXNG3ncv1Z0OEE5wDEIIMUV5nO9VgqIuzp
4aNStvZZdcsor8LGpjlkAvmhLGJzMQDHTQYn1hWxVKOnTp7lvLF8IsoQPBqWH3k0He13HKqBhh6n
GbZX6lgJdSCREBk8JyAFTrQUe3N2tjWYhC24Y9LMY+SQ4jgYs3OwlZp5cB1UF2rk3B4jepfryzP5
Gckg/PqhWbN4oYN4VaocPfB9dFO14OSL1g/rouMHpHgJ2jQZ8GvEV0wyCd8Nvajhu3Df71q+8tMD
SGecNmEKZ1U61GlPY3hmYZeXpk8LmuyY1yacIa3IiUmhcfLdWuUht11PdLGtp00PGRodcvUOcpHz
kk4r/031VACMdjsww35RqeuwgTvSDLjdmVC74u92dXE849+Kj5ND1FzceLs/dlHj+KXViN07XOFx
pfWccjjjsW8/PDkpNvKBEdMnXDWkN+yI2LCgDDOfgSDE5jVjynmIrXsLPYjyJDv7SOxVx8hecjF4
YqTjfeRC95zPxupRQw9vX0gO7T7b9P3zZ1OP7PBN+DOxyQXUQCdWVrAmUA+LhSiP3geOq8ELsadx
qlb7KPIgTAvFZcl1StfkvvM4viVZIp6ZR5A0AANCEzxIc8DDGp5D1bKQslmkljWKR3+ovYjHaVsO
Zm19CRFmroAtKHoZ/EZfhcZhMfFZm2+iqUu/VeF74eX1rs8WNBpKa7zEbh/BOlBIE1Sj1sH3W1yR
40OZs5chfboFXkgJEW7vrKxxLILoMP2gTxqKZozZ1D1OBncVWmYDx9HpRI/Zvk8xrbax824r84Ri
MlQi43nJk3ikYaTB5bzpA/gAsGpZCOTk/+ozRB94KSrDOw1YLDWbI4HyK3suPuId7x52wxsJ/yAR
wSgaC+FqSvvLLDtI1ehMoa63ndWM5HyYvul7DN5PN/mbtYc/G8uQPJ2dMF9j0ugZaRSTrD58IRtk
OsbGfdV/zuq1q+4CiYTft2qKoP8lk/DuRxsGDZaHum12OiNHhTJPHS0M99y3n1hI/E5RXRhyrKtB
oHljN6JlTd6c2170w5jVpnKMlOuSNe7w+FWTd1mgpsVNdkLy19gbeiBh3dt3N+U5ogSIkRm/e8+J
KMBKjkwF21O2DnJl9KwdP4X/NSvnGkKCISMJe7ImQOVkfIqwX07DlPT2t0X0hSUjBkyCFP6K9EJv
ohxSBxMLu192RmZGDq6o1uTlGDEriwxmsCUHY92a+p7WZpUCfGyy7/cRX0a57AcF957LqAYKW05p
VD3w+UfLLCdmf1MmsveSvN0Gm92iFkRdXt0f2T8lDT7MTxjAv15XvhC5K2hjFhrD1q4KQpKfixAs
GgPaebrUWSPYAqnRfUyOSOCo26NWQ8vOkdyoAR5+9w7M3Yyir7EznX1eILqjHkeLCUy//D7AhNz3
Nxz+m8Mh5GWvpNM+/BqxM6AfTIjT9OwWKYHCJj2rqvhepKiJOQ8gq8v9TAoKbvO429Pi7shdcBjw
92gJ3Q1LHohqUa113C9Y6EAIBr7DvDqAcEghZa+a+SJi58onIDfJtxyv/DrOabAVBzNYSoTuTeQQ
Mm+E48SkeyY0/dYmR0yUl01NOzkbTYrk6vu1VfPZ6dRjNHi3opGmFRhSSutOqCLEkSzh6Owj/mtI
RYAnWwfc3MegKaBs6BVxQ4HetEmrvGl4idrysOwfaL5FCnBnmLCfDAhDNFZ0Jrs3r4gJjtH7IKhD
C8/bB3JNV/TryYGToAffuBVmXZLVA6keuKzqbLyOz5hwJA6SVxWn6rbv5kkHFomG6bXNV3sYUqg7
gM6SIeBUdHP19fzkJRIyPIGHkpdthUoqMbtbH+UAzbEPi6rKRwWsmbRgTI7Glo0UNUSDbPi1Fdmt
oB0l/MyyxZlfZWmGhBeEfM4NpT369vCD4QEZcXH0LluWUGYGZmiislfoIF928xVbc3C95SGIkjA7
3lFMSaV9V3gA/3VMs6Phl2MlffO3pEibWmHaioGWaVhZBqskauKxHqwo+3sUgZICf0KLwNkcVZah
fnpk5f08QUCCHfdFCisbzJOfchQSEVs4MS0Sbk96quXUe+/2FVcN1NGFweU7r6xJ5WCPQ/6aERdC
SWJYtF9V6JFILBkkPPD2wEAR+cgg55XJEbZm1jkvrBGoxMbICkhq+/TfNf0jGHvXogzBzUe6aRLd
4ZUezKehP/8fQXIWjCRXfrPYZsTYmWrU9IO63AX1kVcri9KObOEB2/GdWkSkRbz+OwrHXKbKA7xk
Dyc19SKc4USnL7xc7pMhuG5g1uLols+TQTHnkwT4FH5i8kyjiiiTOsY7W+AGZHUKOiTTFCGxE2mF
umghpRo5Otk7WXEnRAZwhU0hPnjxV4L2FHErzQmQrzOcdQwiFoVKGLvuuQzZ9T01n3udETBOajyX
vq5uAd3TTDbnMvbSpsM+hFbRL6FkXqguBaQSD/zbvHlgshcnAvUc6u6m2zlmfI5GV6RH1FqP+i5T
vltqaO8zS4ItIv0dTKg+Nw1SmiiaTE5A+0EGwtz3MOo2UQ+8S0JA08pKktaw1eKIEtLp0FrZAE77
GG4J1sT8g0MSlOsre4eRpF9C+DMpMVNRctuegGtg8MwAav//ThlU5WQWh3mCCR0JgvaHvT3lszaw
MYMkZHRtduU+aw0gBunW5H6Ypo8isrV3TmmokH4qvaTbQ9FuL+q/rP8oBDiCXmxS8txsVKdMz4Ks
EMNk1khBuNnXHAo9Vqj25tPxd3I6Ea6/xxqIgw23bPVTuCYp+CfTnzBhHJM02zK9iyrQu9ltjynd
kK7XXIdDrdtAl84Qr+a2RYHruqfmwTIvnMaJIoeWiAkbI+cs0fd1ez69ol8azgarjkO7vYJDXpUi
yo7SpkzlIUZQLDtmJpS1NmnFGJb75IVmwO2DOFS2xheAfYHCP3XxkURlHDa3QNkdpB0bLjk/1j/N
jz5cCJgQY4kDpnFepTTo72gNdYvSAKr+AKwYfr2NAeBh9PV8NYDHvg7rEXT1J6WhRa/ymjyvfhU7
BhR3sesEDi+5obXS4TtMBRwCUEf7P5BuOg1xiDYpoaWRE2NZVAQjiZIXOeJtBY9GTGYf8SswxEsp
oXSCx18uh/oieU9trGjM0WVhixVqlm0Rn8lLBmsOAVpqtqGGh5Ef71T6YRVOkZGpEOKQSDUjhpW+
A5F2+MC3noJBCoDRN5IHK8hc4SqobofZlN8o45GbYHdAiRHMzM6b0eDfV+njdaWxsi/ePxcOVIAV
SjttfIyUzdVs5cv4HE5Z0TaZFACoppz4UJDmzl3PvrT4pwtuQhoCJj6B/5VZW11/4IcjrGpgO1fN
Wc8GPpQfyLUScloqt9nTAf4TkaSL9tbPpFiBu6HKKKThB/5unAJR6YvyxgnxuZiGuMq3cdRUZDv4
Jb7JKyFjiXAhr1CrXLcJ8nsoLuTviqD3Wj4S0swlwZ1PwcYewhIAw2kV3Z3CRF/PkZEuRAe/1BHm
57RxW+GdK1zmprlLJu+Gjv/lconqYUAFnUb8IREfB/TI+Z9QxOg79tG68r6KyMjAL6q5Eew9sipy
b2cGKxG8bDkfLXJ4lOSzmaisW1QuJNqHBqOR816kZSnEUQwN+LkQcEzq4wzcAtxlttbtZGNhAONX
lr24ZGW375Ya1vam96nMzIxEf5E+8o378sjNAPzkPKyunfVX7fUGQ17KU6T55CVzS77mKAXxiaj6
pw3cLE/TzPBuGjYI4mEEjIxKY8fOfZkq9gVCWGu7Cm1IacdZKpDXBLUxUBOBI5wa6mP1KlQ9aUR4
w+19MiKpw/n6MU7sKmQfWNcbxwoTibw6AkmRcq7kw+xc0ESB62TCa+4+YgdZq6gjjeF12h43ymfX
RhC5wMK0vy+0plKQdGx8JgYQOwUoCpJeMs57W133tbV4ojwTAg8ULWWBStv7ZhNkb02CjF55CBlO
8rzOh/XqUF7sB7+ZdNa1z7aQKb75jgYYsd5rKQDkZ+Ie6KOERfHL3e9dOEaNBQr/kJPYBPs5bavk
KdojInZZKVxhxHR0wFsKzx7Qb+Z8LjoAEWRFnMv+vRyx+lkx/5e8/GfyYuMVQXj0pLant2VFLebT
/6MKRnghzTcB/8808M22+AhrxeVxRwpPvxWi/85Q+QWRYRky+LkdlOq2YRpkxLVRCNsim3pwkSrr
BAQw9FQEIyCVQ7NFlKbon876Ndh/jBYcodIpFCzRK5tVtOPlwetcNcDOSzb68RUEUbFk79WY52/3
OA5tfEv1rPyAn5hsuw0SMAreI56YyqtzbgqdAb0WMrCys8aGWILjOuBLSX1vo00BVkzQC+eFZhAc
d9KaQk865Xujnl2drQhOlaCrCYzNjivRiGbEayHk+2+CS1KlAyawOX2wpfXl4XXJrK8HyvpGZ+rO
ZzAvkWGdehpC3nj59nWTAVV5sXOI/zRlYdss9AX7Myew+Y4Dj3ldeMf+nHgkyj5qYzkxK164XKFf
VCZ8hoteTu6u62bBNtAQRDjfCZgGbzPWCaPM1G0dioeu4MskOHJa4tIRfr995+nYCZH57QPKbUCq
0w6MrZjMkSymee3Di6ar4fZ44q7OYpwNOwlH8jdj0YKsuCLJHzoW95QCLEbN2PGTZKUA3egU12l6
ZprTVoA5Kjjr54aHJu57I1sAutVRw40rVQRax+np9e6XclfBLAy4bVop8VaW7SsXhVJwnmGTrAhF
T2OA0510C/y2XUFIQ3D3pCqpTfaw93OgxCAB7bqm78Gq5P/FN5gtRzQd9ddhVZZc8Bl9Qdf3wEuf
XxgB9NhrfMe0E38v1OKQMfpRlOAfcyX5oHSOJuFWQ7+FCmAAAggcMN9m0GU4xGV3BL4FXpNv9ruv
/n+HGzkLxPTFm7rxG+F5VLuPBRRB1w5BZi2BoGtwxJej2PVjvhIogclJPnqwx00K9WWudmiCkBNR
YtyU5sN+FklEpOkWFIn6/U99LE7CCwGj42oOnq/zbZlDKuN9anSKFStFKs3VzL267Vf8hLFWp6m8
FN9eB7mZLXtjUoYKayiADYQnKRK1FnHtxvA5W661tafYDGCt1YVCnrANLf8q5mhcuxnx4TJy3zHv
08r78tPWF602EHBE9U36VtpdhRCPvkPQUFk8LUtq55xdDnKArQ15N4iGFo5kl34DPqOtKeRdVMwe
TRZNouVEuaQVvI31JpDsEtsiTeLEvPR3tfnnp0yNeLpKoDyZSyYsoG4Z1USLcNZ0cz1sQdfvbr6h
VD8h1rzsu6NYJZjdZb5yCTZWxETbQoxYpRCjjzFrw0/Jpe7xT8jcoPNXqWECKBufSELTGSwUZXMf
a0U5ksGV9O7iP8f9W+jLmgLq9IHRvv4mhXoNIi34uUi+sqNwZjC4p0ZFDDg2vEmwGqI9cCq3lJM8
96TV/F4huO76iubYuubCfwWKRZDLjnUSe68W9dY4v3NVqQf9Yp2fixbH1xNw5nCQqhHpgY6KIpKj
Bkbl2UljxMalqtYIR4poSsK/Mhigjvy6iztZXIFGStAR5FUbyD2omhUoAw5lEQIiFelH/d6w6skt
cUZJgfNKMEUErsUGIi3bRrTAxql9AdPYUQsEPHROWdrUGNlAOhIlnQ/O5aJ0psusOJYnx7db9c65
DFRmCrOFX35ndyTqFVvXOpf5acthcQ44n7qXXp4dxQm7fms64MvarSIb6tSFaF1TTVHsngyzXoVZ
r92OaAvTvO0s9dBZ0A/ukac65qZxQfpqJwspHgpUcdwCGPQuq11FD+1uUZT4eJAd4DkjHHcIYGG7
97KQQ1btGGoLEqNjgT++qFqsuv3J1HrlqCcQvcBcYPzsRrRo9h030ZVLAirPBZHfX7NSOt2luatD
Pfjb0NV8QtDaFjieyqOqPu+py9lpgN1zJqB5hn1/uV1AgPtkvAmR9chHcy/352GgWSJQSwCPvKDn
WzxrMT91nfOP7FPMTk0za1giyPb/f6oh8mhz/MmvBmu+olv1N7Dd+Cci5GrNZh+Iz2dRWGqSRSJH
pIizBJD1nHzKgVXsyYc6Xo2sJqpbyuR+J7YSMZrtTOMjlhQUKax3H+gDBNB/J3S1Bcg4Rzccu+2s
up/yM/N2utZVcNzyoWVBoxR0aXifVyBnd6X4pi0WttCqJp00opueCvVusfg2gbycpKSXlEdDKR5T
D6GHBqR8t8+rQIppzFrnSVEZ9SK9yQEU0oCmu+1tDxxYUjbZ50mbHZiAGp3H74S9GpqSNjVj01Gu
qsuB/rl1B1G6MpR0tNFb89fE6eo+MuTDzSoW1Xfq6iI/OCCnJsoZeoV7aSvo7KD2fTiHWqtQkYcw
FCwTxxag2yWB59s7Q3V/5q3AAHAop2cx2Dvdwb/MvQpXwwuGHA+Ca/LruziQrnN6cRUAp7hqFp0e
wPb7gP5o73fakbgm1zw5aykW+KxYri6yLNohr1Rj0YTI5cwchuc0fYbJKeSCuxMyAk/3xOSZuDzp
CCu6RL+wh1KRyb7KsaHmOTVQHD6+JuiYskOjtG4wTrXaYIUhDBelMa3ubiIzLGf3uFCGZjd9Z63C
RypJgpwXIEgGhE30eeINmlI5sKtZCW8nGqS6EWb2rIiiIcoOj+AnX78QP52WAoW1XoNb24FkNTQZ
UWu/QaUPsXlNaW8V2iA3q+RYkg86pSwsbuDFBHeBNGJwW0m0jZVUiUvhzQtTvJcZtPp3cbsLCmMk
GrxqEWL224zsXic61jiAIAUg6/ODlezTAeH5VWIfAFGb+pxKk44WOEEc+X20RoVu+XMaDx7Nrcm8
2p1lU0OYisEOaektR0g5W1ZAXER4PxUXJwmtuMC3v6keDejL1Zq0GeYwD3isjfSqCo3egsIWu0xY
muQfDZG2goDz5OwF7UtJg1wS0St92o+ND5O0/AvcLi41omgAuAocVrTrGSEGtG3EjTi/8x5xSnt1
FCbiRs1oNKm8fA5CAaCgQKJ/8GqR3ozeBUT5xFhHaF7g2G4Xenx85Um0QUdQWEHk5yrYszpAwHNX
Uj27plY/NSjMQfxKtZXnv7ANWwgX+8GlopDjLsYrO/OjRYBbHfySAMYcLnl5sNPxod1Gp2vTUBtU
E6l6fMq2x7RFf+luAe9+xD/w2pqP4O7G3Xw1rdQpU/EJ96W5c+IPCs/0A9oH83YiEU7ZgXsyXfMp
s+xHb9DwxdezFS7Z+Cf43zNPfOal0HynV8oiqRAt+xvO87bzuqYH4c6arCaKUgN1QOOc6fOmPBOa
HviqRU6C2Skkf6tQAgyg0XVl9ct2P0CzC4/TZIb/NVwbkEeeM1lvZ8G7uebL+kIqNpgsK9lRVShu
zyBMaghkKel8Ho/FuxBr6wrIK4KPkEkKIhhcg5FqjLHp8KG9wxmjbYacW3k9hGC3x7y25NGW/GgO
DT2tQ97ufJDQA7AGTSOsF/G+Pxw0bDFasbz7kY8QjsCaoUUTg3BD3aee1Q+hDWCjiiWxwRql4aEe
qodUW3tfTbSkbjOoGhUK6TUlItRG53I9d1z74OFqy92cwfdIBuDTA0BVcHzvJnxi3mdzOwKVhdZS
rQqXFEju3soMWLUO40K/D4gSESqYb4BBqZdb+OnlTXmx/bb+IaMk+mA1RQFc0fHsCy1tDCqP4C/o
2nJN7dUTjiCC38zBfO+UigG0+MUi93Fu6aG6h+Cpf+gEtZiS3rUSysjtL99zjzFfCEB9TycAWH2r
K9Y7/BBED3P6V7+yrzM7JpeAiXLYQMU2Y6Dc7xNVSqaMWDG16Dvit4m1TDnW4KSfVE8+woxpmjrH
XBL1UVgn/LO8LfNICq9wMHGYrj4YUjnsdQK6i/tSIObZxSSzZvLNJ0IJGm/M5h9jTZ+gWl3AQOKl
mOlffBRGs2L0a8oCWYaANgi8g/tx8omQ9PGlYapt9Lw1ZBte+2rq9TPN3QeW7PCaFlmEqLiQJMeK
vHPnn9vsr3bGZInvnOOgeBwBPpysSpWemPl/KPhq1I7e5fFVWpTGrjHnb1aXAIl2ZDP4GLTElJic
5uNq36FzEBOXMCOLAygnIzBBotxiHp9oY4Piczg61/eErPCGjjWWtMcOeT8Al/kzRI+yEiK5AeWu
QZaN2ALo9wDeW9jBBWR6WwXYqGqpmYYJ/9/LiMtB5/ew+F1dZQajFP5Ngllg8dgv2R/+Z6S6Ah/+
K+2Fy9tEGGq9SVYDtFr6fON+Ci8p8LHfU8t8fFMORt+J7yg6WY7UmdqND4G19t4TkLoXmKYgL1Nz
r5Ezxdgcwp30+zqcTATaq9kJVv20YW4u7KFbd4FlFm1UwYpwHdBYojPQxJhKnQ9a74XxrJtmjjgT
PXALQYiN6NaDD0gwm7lq5VhVYWVtjGhDVG3VaZv3eLpdM4ZvWQa4pcEPVz4zADoYjtY04mcRe+V9
xxuTESi8ejTTWw4/lLih0H/AcjN9xOmfh22ZC4j5mzBvA8WHVLYTch7XPNx++QsgceOE85eGuEyq
aK6bE172ls7nqK2YCuv7/Enf1K3WttSMFi92/CYOkCdbu8NsddxKg+bGW13qFRnPMRP2R4N12rZI
rs0mNmJrDwGya8HsqUbNjI8/SyntZsHfANopmWcSOOXv5m064e0cX9Apod/e8bBakw6orA20tsjF
bhkJ2tzWixPIr5QBcbfghPnjPBzzeSsNnuNKpTKYVt0ab8V2ORzvUWgYxcHjBb9B2Q/wmEyXFA/5
DgpeNeQGCTGFoqSRXAGMbfZTETaZ70ZLOdr/iY9zJAvtxGy76yUHNMJz2acSG2s+5S+/EPCLdACt
pqczvPZZUmE3hkr0y4HXL6PElSwkveRd6XdCM07tzTzjeKJfy/ccoiqSIDdVjBo7IEo9DBGcfaGh
8qGdh0HOYna5I+eTAJWkcWA1RHxGL80S9kzXhTEzve/sHX8t7iNXL8JnY4tZiZUIWRX01SMrAnQx
1jSZvTG23jD7jEvgKqyXospEXVxSjeHsP8TL9/RlJwHPXlRaobSy5nPXUYrhNfr/mRFuQLrNanoz
W28cFn2TlPkfZjs6GFgPfxDRH7P9RuFwBviZBw2OtQEznS36KaaRxOraELSIZWNxshFuLa1l6g5v
T1b0ajYW6Hth/SvejZZU8B/ub3x4s+TnrMYV3qM+D8S+YnRFzoefq3Epjj1AoBdvQYYvNxPEI0JK
8t+ha9BSTjQdzC6vqtta8ECwvth8fCAWX4UPjvD1jNT8DG4hZZITUB3kWUKCFwxNxaucMDTNRT6v
Hz/iok/ETK8SISyBp4Rbbdas4i7rR5ddDb8o33lkXQvHUc7+Nn4k250sn+U4dty4GgbfSczwT5xU
U6lp7gCVKXnJjaGa+zR2rYLg/IxyTYhT84Jvd7ULi4ft2+bFw0gSAqJhUfnMNXr3PF7qk3vDcvc2
8OH7G+SyEau+PkUhzPKylQXkSk1BULepqGUyFDEXUdPXYrNSoYPHK7/5pKBtVAZ79b3p9/qusY+t
F2O/vrMUI81GH7mz1d84mu1Z2s9gtTQjMbJzjjs0CihtekEmjSf1lnWmdKavA7PfwA0N+mLpwtqB
g9GkElIWWp0A13ss+vcRv3LBN3WmAD3Zq5OkbA/wlZvS7MEeG761cXYJimdIhLvGJKSN/EUo6TYC
2paztZMM0Vdgd7Raa3tmSjD3v8G9sSq9OXR4piLHXE7ta7xqggofPfp91+yz9HfnbHWtv3oAeuP8
j88eHKozf35xEaD2SruIKT4EI+7e66uFTL7fAqwfmn/7jhMOy+Cj9Tks9iuMUE7g9Pn3EHLWfS2m
skSDhBQzBBpDT/QuQBiL3KET9+x6pJTkgmEsPpivqISiqLYLU+kr7Qazbk9BlIONjbhxBb2VcJ/I
yPgkHef98e2QRR7ZBolNOD7mkjC4RQl75AT0pKpLdCc452r0H2pLX1Bt3ral5ZSczTv4TgoYpO2U
l0OezlqAYQNZ4jpUvbqyIB4fcbPmCCHq5i73k9xCpe0mN4WuJ8Ee1Nd2cmWb/w+KfTBG7TNfvpgA
eHhhJsonUmBbCSruOKsVIN14Oh30QgUswZrcb6Fs3FuAsLbl7dRNS6m9+WSH8BzGAtMuNFRj5zhD
VMjY2Z/2ODr4CNfH+XFTu9qTbr5owYDcIcPWx0h/OOs8gWFji5uG0DLdIoF7wQLWyGA9WnI1WkFR
fSPki9WvN2cO1LhYo4LV+RKyMI+u27wvJJx+kHvGzJgf3yp1u+eT7zhbwegUGrzfMbNKzgPWuuWy
Zz6KgtEVs3Ya61CISOeb60v/oPbnlamZ8k/FkAYd+uMBqL2UOssY+n5OPp6Z5mDazYoOIqrYnOYE
OKK5OiFHHLrzLlIkoz815aQq9Q/rpJg4CfTUWin3eu+914lDFdw3j+b1V0nWZ/HpnFM0ICS288Dq
B2LzI8g8YrViRSr8HDI7rO9+9oxWe22JG2gjvX60Off2fDGZzc8o+bk36kGVTcz64UVBts8JXoR4
tMtf9UDtKsOzPtNAuSBJytMzNJHf4Sij62JRjleSChlW8jBR16oMHUbgtd+2HtNU+E4C/fpbbMKd
ekYAYCZAQ+mkJl1e4TKmzSFyM9uuH/RtJylapcY+D3/lrtPsQ9s5g8AqjHlw9ZF9JAN88lQeL/bh
GxyhyZ2n25dx8T0nXuvPmTRlo/3w1Tm8NXlMh/bnpHg72aGn8pBDy/uWAoJZhx8m4XMe6wjeJ9dV
J1hhxhOcTWW/V1tCJIBLifeQmJ5bKnJjPAsg9DbVs4L9lDtGhc8RJwIJfY05lrwZfVUmjs+0sTy+
Nzu9VirwahvB3ZNOwsZQAY79LvFZa8kX+zm5l6j77/v5pijq2SfMnemByGEaYA2ffBeHtllqxlg5
CTUDgP1C+kDT9SiBQsOVI91rvHxftWE2xdSyRq+ej0yhnN8VJD7CoNIv7geaIOMeFV3XgYb73VzR
4MIRa3EwannJh3YfDLz0pbnoQHVzl83QgwefSDlU8hAzkjXJpVbINHxZTEdaVDWrbj7L+NVVMgQM
uYUxZXKaOCN4DUqQA2kZKqVR8cQX06bQb3WAaF33us1+ZKVkQyGgCwVvMLIbRTPOtq8fY0O5ji4G
tjFJpWGx6JOUdYkSo9iucIOUjgqDyiLIOxyGMkfk5/47EhEn/krOC8P9FF5Mwq5W9/knGL/QYq8c
Y1vDwnYXDAU+e+ewZ7vltv4mr19KFuGmikCnj+MZ+j6C9o5gr+2xQLFCHjqP0suJB/9kEB97mXwz
VhpxRaLiL59jkSjHJSY5EZLSQai9owjiZRgmbfMbXMwZibAlDrXaW07eBQ99fAEaDTVIgLIzo+0J
P+6n0Qk1+/3nFENxxLUPmSnsyw2NukPfcnKRESey1+Hiq0OGpZ7pVYxduiutmcjrwNtK1DSOpGTa
yKTNh5GuSa+KdXsPYl9YcUh1SgkQy2Z72GIt9leREIf1C2CUTp5MHtntotIgzkWDIfoIGbf5Iulo
B0s0EhG656Z/PbojUxq+9x7Lbbzcyl6z5lF9i1yMQkxm86CheIp6lQKO5n/cUesefwi8wIUvvhpL
vmREwnDuMbudx6bjumgj3hipFTV/kmXg5iyFeM7nfSA8T3kowMKC4zIcZ13PTaHx+J/VQdBMFG61
eWKyMXuB/WldmovHyp5NAI/siYXlrwcnVv9guJF0Wpam81K0AdGWUA9wjQmG3G5iTqr1uT3pWmDL
QIb0ySL7r+edtHxBhAfMLlJyY1g87Se0eOLfoibMm6x02TvFFJS+CgDnsJMDwiMWOVIR60Y1WHQX
65QfzXjIeabuhPiIgIaF7K6P/NJvn0nIERvIDEwJnNZrVme28o3VUQCwAYCbYyRKrkjvl3LBlERq
A/UPeSzildH/TGQswDGJT/uBNwY1b3QnX0yyqIF1/mgr6xkDapcB4vaBJUwtVhO93mSrZ7P3AfrR
a8lynU1UqGW0j3ODGJ8/2nZ4KZhvEP8RbrTOsooIfpsy9tjzRItZ3rqXr6XkaClF0Z6f3E3+NRm+
OLeAngGdQpqGh3pRzjfWRaSIOs7cVfcecSEA3SDLceouFsmxxWdfg9C5NotC0qzqaOAoy2dB0jKu
tHCSjQWZHaZpsSIdZo7Mg9Ltiw2cBxpIggu75nA2R2TKfC2ErMXWGJL2/m1Otog8xyT0INRIxKsm
tsZ8MDkRKTfBFjfROdDUl0taA5V1QQHQhNF1f7iJvD4hGBF0rGEOYaD+BjLt7N8M/P8Z4VBMne7O
z+WXzJ9H5xnHXamZvYQrMiuMWmYaL4QOLzH13Y8xAZDG9G43jTp0vPxbRviXaJ1mUzGrzgVPE+/C
iY4YzFSjMEtfmO2wXh46Wi1VT9qUKbcgwFqGG+JYiCZzaV4Eghtc2lCLd0ay2Kx+pfanXXIB4pOS
8L7aTduR7h6Xdf+t4NIjfQizClgY61tggdX8hr948Eb4yh+9Q9HUd6Hp8fFjSVcrKBZOESyQBnhE
3WFATVA5W60kKaJvgafmAEFbLcdtWt1XkmLZdprQXO3rCa6+Yyaf9iZZ4pcfjrhJUpMBoqOL7dmn
ZKsCImXCrNBZCKFtjM+CZ61j519AJmcKiZZ9T/khgYAsfAhvgXEqFxJQJ2E7Ohff6v3CjOW7he57
HVGg+AxJFRIg6firQJvkZa2ZPYsEDFxpZBQHPmoFcn5MlB2oKUD2SIRw1ghFWjNW9C73x56+nDDA
UfZ9CAskyF+TrcXAv43CXJBnU9Lo7aT5fe4Jk1XwuvC7u3doLe+/rbgUidweS6lBNUZZfUiLPWAK
elZXUwitQckyaLwlUifTT9DDCTnL3/pXpJjwUd8I7oXGKZHJjvVOmHbixXPkAF6TF+Df23CUBGaN
33gsgzy9pXudPWe7DI/GIYrXu/Zk1ZfapivX/EbaUk6YXLMlHOvXPMopMvje3hkQu1MIXVvKuFrH
+VFKsLTDxFuVe8fXpDwZWp5o6c5xD5bUriqEA2qU+XVMOkDV8Ne/Tcu0y8yKjsSlOHYieRLkh4MF
/mg0Lo4PlA4YqxV1sddrp0paKB91hQQ/srwnkn9YwvccqA39nBCy4Pp/BhuFUn/xCK5E9oJ4toTS
Ii+YdfjWNkWTNGDmXkf5x6g+ApMXGjNtHL+JUSmWU+zDqSgsC5y+hIORbEdx595P2LkvabdK1h0l
WLl5Un+gNAXH+pQfCG1pThgS2BezGTNa1SFF5p2+3FXGxqYkNoKG7BsoYbY0rnsf5gGHUT7TS0I0
FWOhL9sIkP8QSbKn6TrbR6illap0lYFyHYJQ2UBdEXBO4q+ji9Usq8xe/XZyTuuHNNmMAXxuYKlW
IeSms/jXcO/25FRBaXutmJFU1MMdcX5gg5a/ETA3iQC9w2XggqEfUWFO8/Smp44c35qLperCQoq4
zDr/DtDebOAFn7Apnh0YluSC+DVzA8YrcpANJ0qvTKRvmdYFm+gCtf2CoJOj52cad2DRsMUdtCCn
fo/8T2iI9pU5ReFhMWgv+H/tpgCB+cxbre4fJgYaxaLvVOLXa2UpjGIP24AvB+iNmzq46eruzrkd
U1+tAg8+fsWVDeUBSryYtt86XDWfdsoORkLeg1l1f+JSEwmPvPq5v8GwUr2Xc8K2/0tSRCXg4emz
jGmHz4/cpGCqu2OCNe2n7jK4z/i+KWG5oBfVClBbq+BndOS5BaAZzAz1my98DT4i27IrpvytsfiV
lihFUo8I2eEJA1q7kQfmfUP+rGNxFh0mCC1RDyS9WcV/mpHRZ6nEQc6g705bW1iPT5EZcuEunLiI
2LICPSgFf3xdiST5cRkAwy2FralfIMy7asaDD2zJ2QRgeQwx6T8lJWKC5DcnRsxvU+OZ9OWBbQKQ
akS7/P2+4hJ02XGQ/rXoRGoKFIUlUpTRas1QdNa7bRGVftfG59wUzNCeKj2lR/IuUVili5C14OGo
7RcsJWJ9IrGWajVYZRn1wbECT38viNfUTaTQ1azXmw4eYZTsaNCYKXe1Ku9wZupmOWfSQ1jkfMXa
mSyta+0hj1+dx1oCPuAz8o3xbM0icWydPxhPgcjppCuTvMfPhLBS/ecSaqoB1nto1yr7IKH6BWO9
bKJnp6Yy6lHPHK/bdd8pvs0ptKm/ICUTVur2kC5fbfBiXqgn4ezEaKCizggZDY4SqPoFB3Tdbk97
3ErJDH2gFDVjHA+4eGsnbw9wmCIfWREdICt7TV7tEMYvq2a7VM74z4L4wOVDFsVvAVTCRAUSiKu9
Pd3rE6npH5ukW+oypXgTSPXGRR0liQUXVpDqf5MAJuFoIoI5W5efOt1s6Fuy7qC/8oTQP7xkPomC
fuXbwyA+j8J9yIvBXDdhv8brR/ukKVPCI/02+asKuZePVEJHpE9WDEudC6/UVKbpYBvMkzmRJE/c
5z0IqQ74BxeFRtwtjFksjSm13iKJSDtGCI7fNThD5NpG9IajtjwooAt2z55RDotJOTI7AeIe1m7x
fdlgIxyWDVYn+23q645mASFLBN9pzyHEgOvsgOCSQCsPIOiNtFiFQ0hcGvrtykX9uqZjpaueppa0
YecxcGnPPy9m3JV7zcGaxHSOjYeqzgio4iLYefpQoKF83eBkTK7seLI2UfBNB6k1DV+deYP631na
Fd7XM1//8EpdBWlad8GIK5Zv3M71McT032/KhOR+mlAyJc7lJGmGpB3maIuw0tqjdtTAWqJt0klP
eHZrrBSfJe+Uezqqw/ZE/LpuHE6y+W41rxwBgDJ1uRkNmYIvqizQDgHOm8xoS3i9YH1gPUrBR6pc
kWKAsx1yfhjPwQiDbGJRRhXbpHiRiI8w424OHOlsQAOhkrFZXaWgbOo1IeAQE/GZd7Yz90igu7uZ
h4hs4yd4GKyss4wCqbnlWMKyN/aAamv/p9xB59QXQpTNMYZlMpq/bmG9KCeetUDuKsAVZdoeTLua
ltqGyj0WIS4LIbjVrI22o6BMSRtTqkgiY9wuu3U1Fcq3Z5Su4aPEHhaNaZVqojBiGOEgRkEtIB6U
kU3Sw97KAGnc4hHZg45UkQLOzZuN1qQ8n1aNjpSu/btf/8OpgXoK9heeSi3z/LaUZ1dEcfxmE642
3+hDtrrYZPchZAV4CUm2tVfYDI86TYPoaikrmA0w0Nt5BX27aoy//P9lVp82YUZ551uYZvMKo+hZ
FSOF/PofwBhHUtmQdk7k9BabS/vnIECV1J7614WHd9H/uuxjBmtDr8+z4aUO63rfUc1MlaGcHdxL
vb2jPMc9kp8mQsIT1QGP5v3jn32v0fkByVB2esPFNLOVcuZD4scgcSdGMGUpsezWIDdI0DDY5Xah
O5sgAS79xfvujVBlDh/poYKDBTUagIj2+yYL1HW5kY2//VXZ0Mu9VP2LdIcrMH+SoCmOXp4ZlvvA
dkTO/0OZSg6s/US59lYTkDgzs+oMb3e3raa1BfBVLrPCpAo/DCKvyvvMmgZ0/fXhBtLT3U9rqoDp
VVsTK2SygstiZ93fJukJ0vJdvB7q7+ZabRR2uT7Y+hhjBi8Z2w+GBgkOZQ8eUI+6dBeUVnx7utpf
8Nm3KWCVJXY8IKRFOJP/KRmaSB2GIiCcDEx+Fawz88mi1zAz5PHImatvWfTfRaCQQ4E7Zrz632Zc
446AQm6nDs2SlobEtrXuLUB1iSYWo19FNQGpQgmGi+cazVTwGqSsTimAL+M5PwugnJM/dG7YO4i1
AARn+1eQUjmRmmbTgGgiT/6pKXlvKtsf0nnf4bd5KX4jifuNOiBDy0AmXxEbclQJsy62DlFxRsiZ
yNrjbXWrM8GxtU6RNgjnXLc+1Asu8SaHSxyzoJB3//WoHq8aWLNFtm8Kv7YG4uFd3PumMVBbPZTG
fwf+mcGOFNEVAuwGVacyobMqroUcZgQ1cEm1D8l/YxnQ3xwsNlKtwOmNSf3NdhQFaJxWgXQvfVGA
+igYQnH0OunGxrWLnmX5NlpbZWDcXhizLJYVME1B5bD8YPT0WJEr5CYJTjg/33/0k9AmAqR8QdqV
/uFcK6JNSHQ6u3DMQXVnsYU9QtBSl4csAattLob2R6Ck5JT1oSbvji/TKqmASWf0XQhLHrvohi7e
rKtbhac83R1nKFkyBbf728GnSfoyOTFKLHFkUjno2gWIcpcY0tcPZ6Hz3KSOEDXEV9W4XAZoST24
2poyRc6655+xcYWVRnCkiY+FODkunzlCpo/hVDXZgzNaqkdmos38rsRKQTCj3YXm1d2DN/NhD+4a
0DPGV2azve1Y1NU41PsocLbVvoUCHUNtIuegpK/yHLSGmUP8OF7MHPX/RLWDYdOdOfP6lRE7vllK
NW01aoWCgrqtVoAp3LSXK469mlzEaSdqkOIgVAyd31meY2N72LU8l3Wqd46TeGZ3YO0fFmYAUQye
m2WtOvSIo6BXWQMCpapwuLewaN3cj62yKXNR0vANb0DnkW2NaKwmKC/5sI/1xOb9ZuBHdvgRBW8G
+/DggFft0geSP7n7yWUl9hYIxd3kaBkyPeJsYK7clsABYsQYzvkEuEYwuQujH5tHiQMbpMhcxqkq
BatlwrjysUMTtVl6FBKmAfgLXieGWdTQP9u47Q0cV9rmiWtUH09dTE1yqU++kulOtnoMNj6woJ0F
4M+hEN4A5xN7bOQEONn4Ol+SLKVRcsXfg8o5oVN5ch5StpA7iLbG/t0BhEm9QyoiOPfxAkP7yo1f
d7Zc3KGmKHh0+bAmmlHyegA1IeQqNMfP+Yt81PscRWf/kKmXKRh7wnpyDKI3C2QRDUUaTccFP+6V
gEP4qkrSOWhV0JBrMnHTsI1T2Lkbxi99LGvdluJxBkev0i2mkUYjmwMe4xIvzxWMy7eh6s98s25i
/8lhz7bvfi0FgfxkUi/vg87F5ePwOXq4NBlKdCh9IWfCJHpRdPJNJgJaszRi5Erc26ZiX55d1ecr
urRCHaOUu0C9uztSg5p7MjSC+ehYl+ynVg/QatN9uL6SA9ArysgvI37tdWN2udp2zZ/gAw9HNBLN
9syedykHfFzsxPARtVuXJMynoMKbzULpAfMMWUWRHu8MFXk/GejyCcGFzVagaTBLFPaQx5QCYamW
VRF6w0lPNDipNGAiLcsHTYqQ0plFOFEF3thDdAUaKUMHBlGMlDPpvILNeuVWLFwgfuYkp+vG7hHq
LQKD0ehhEeCuPuwihe4EvUYa3NKTnfjIJ1Qmb0rYNwqIy3lf+7+EStlsYew0FT8r3egkUxiRzi0/
lXS3YGOOW/IAqq2pkm1LFEk+UHrDqJNz4I0te2FkWJFwhGyLz65eZ4I71060oxolgthIofEUW7Wb
buFYrF5jmCGUyZ0LYlnjnA9R1rw57e6Nqi4neGIdhYCH6hnW+7dFyCFFYg8zdMHz8UcM59/5IkGS
8HA9P56neBn7XQQTBzN6Vs/Z5rXUNOpppIwU1Y2fbymPkdjsRo/by0xfTWDVLffE9fCPXk2uS+1M
VjFkrPq+XpxiHmTuOj86fDt7pLv5T3hikk1ZxCx8LXeB4SxSjGQdvwAEIQjXypilgl1HKyIQ8zLE
1/dWKx4N+CIGxwP4cLzcbgLSQePuRbK4THkPDcrJZ3GOJBODrseNyVVCL0qhZMn8A0DavM/Sp7Sr
BpexeitQybYFASrTBeEzWPKz1wXg7vr+/8NM7DkI2iOGspmok7zRpVkE1oQFVougRXSieqGoIpcL
qwBDejpSo4fRxGMlBdcuEa6DJnSHVtdsvrw9Ls9lXQI8eZ9uBeNwztC/jhPd3QqyaSq7O06+3OR8
r85xzHNyQY2ey9hSiW57QbSs35Wly7NbAAND41zXk0adIpm9iw6Dkemacq6tsepFxOO2QdvRoXnz
GaGtwKWeJNM2EK7+HxACinT5VrxUTVM/MGjAuBNL3G4+yAj3G5ZQFYU+CGnH0sv4Ulu0+UGy/l1n
L6vEw5SM5vekkyeVBCyexXSeXpxvE2bWGaou+2oxtnf/KTteE4HgQlQ7zxwrZXoPkoNd81YUWNDj
QVUlczz1I7w8rkvXYi0SOk4myOLvC3tTV9ImMQk7Em/gwP/dBw8kkSpeHTHZvshc+5JH7TPwwsWb
n98Ee1JJIfcTeu/dCEke0NQPS3SSn39GfI4vtbOXwz/tTfZGllEolDYR/3CSV9pwXIfwee7yAG0E
Zrv4On/E9V7ZJWhS0WygxRFLGAGfWVGITWgEw7Zc/8x5Ab1/oJ0G5ovfloiXfikYhe61cyggECFz
fDCM8+PNCNsYmf/NJO8F3nwTk03IfDTH0Ae55wap3FVLmBVLnqaik5B4VqBWAgM2GZ2FmVwzmcvE
XUSPRNQkyA8TQGqiFiED+qZSh4iftVcG46A1PjKT1k5Ys8tZYDqdctP9RW5ZwEh9ESLtMRSZSo+S
P60Loj55ryupZA0klku6tBGNVKEGoPDbY7bNSwwfIiNPVJDxh9yNjb5QkmBi5W3iJkCm/czsC73J
xv8aBeehRwV/xEtSeASiJnZGoNp8a+TY4K3slolKSNZYbEN4unNXEQM7BLnsbdSg+hVMqwPdYalS
3ODFuanyh5E5pYF38dLXgSzEiNNl7TbN/pmEsoNQg0nxeU9k/UuvZRd3MLsTRc23AD0CrxRw9tUi
qaO3FZd+8V6/T++90piWLANMmg39aEDrPomt2kSYRS/igcHKdUCTXiGoPWtqAWjAWD2aQbhv6jrK
xFmeSKMIWBMhdSGgY+ADUpcSHXTgUYMO3wnEYcmoWyGXll9Ubfc1uE4SsIFfWlhknUtCdynxAipY
D/fE6rCvOaXpieDtGmPii+7Gty2VdTrnDlvmOUBtY+vL5gJTjenQcK2BC5gE2bNkFGiS3I+pvDZm
WWfLgb2PjrsDhfcmsrCOrOkHiV0necETDBKZh+BwUd/5rxPC4Gc5j99nPHTN3w/VPxXaZqjr9h+w
Oz2jtHMrIfJYuYD4z64pONR99jk3hi8hTPN2cPRCB/3PDmMHCE8rXBlbGxk+hVBEb0GWlU57E8Ji
z/srsLzh/Tpa4A0JkRyFinc+72HOz7W6yUk06Cc4BCSGQ7CQvtFOWaEBTLNsj+ksPG5qhV3Jf0aA
tyIHXHcytYOZoJOWUUXZego2D2so/DBgCDZ3UfyFJjGddZYARXf7fn6ckr+usxjyitbMPIk+IYy6
oA0LCi1rDo9KjtRKpOBODkqtzfnXeiC26nP+hhhdavf8MdMt+xjnBSbUlpuGRfpN9rk+cou6LmY/
JMoO6I0YSDMxTlzJMDidmLbggluKlyopMebV5nHIbwLVuRLRd3h/wVXg9fbk4SPLCmc712kKxd18
mWE/8/hj8zVzUu84Tlh4okC0zLcGcAFfyIxFekKMQfrF3NJcM1TC/3VQtPWgWv4Syj+hgt1zCIlS
MEsPP/EOvvc0Ab+N39JV2oC0rcm0fs+OKBFfg/ZG1T+vM4uMTnAZ1/DJAj92k58fTZ4S+T4YNvuu
bsS+jwWHe3ye0ZBPDyenpEdLxodJY6hc66gVyub+Krn1U/1HpYGt9Eix1jdpYTEt0C4QIhlmxC8/
dWvtXxZ5i3cdA6ExXJkXCpWHN3oyisOnJsRdAShJVvvAH44VDs7Ffy+7LgfMpSy6vBd18OgYpdAu
GdY+qjIJD2Q9TQOpx/1Zr/9vTh0vudn3E0Yrqd80xjDX8Zy6jd1hh8ClMbMUZG9POW+98vqUm4KT
t8wYzLfE2wrWrDwNG6yNrlCkbCaLuHPzByvxVhsIeK++wjIPRnn6CX7d2GjH22YbkfUyqFAiaBFA
stR7kX0MAVtmtIQfoXF87mMbY5OXtwAuo5xMY6ChjjZ/HpYN9yxKdab/R7Q+edXSMiCfmgOYERAH
8zTp9f29oZ9yrXY++Z45xOAq5HFqeln/YFT055CMLeohPJy0ix40KBGDNL1Kc+J4azbR/lHNKldx
H2hSnDC7s8CygTKA5rPkZdpLdxPocgOelyaG84kOr5hR7JIYEB9tBNFqgSmNhx+/gZ5tL57d1Qqq
C5xL3VD7UV5KASRVK35uoU77nkkN2GSxtaZkOcZ3dBNZ0BID/pqCqcUrETTSXstmx5nRSBG17gYx
gsND3QExV5e15l35pHtXuWLvlp4ArBD3ayQP8+u1AnIDCR5Jda/3LXilUm+iR2WeMpfOkM/0QcsD
0i5kMt5OlUvXFDnUuQpy9gN3LdxZEkYB8byz+Af4inhqmdjpbZ0NJUinKxBNlVkkrnR2E9oXho2U
olchlF1kmjj0PvxZMozlnpk0OgY5DhQK5dHpVgII9UIiLfMR4ZJSizj4uKHmBGnOetqv5uOlzgpG
TAsvs50K01InzszLRpnk0Vn4kXGxkCfBBPJrhDw1BcOK50uWZpZNyW+iOkIpHhuw75ZbXhXxXBfP
FDUr9vmO658bPPbP1jJSs/muyagT0phw54a4R0osxCAed0UYtnbUzLh7uNRXxNi90Pqv76vRKNOz
hmxFZkKhyxIsAyEKLD2rV/X6BUxmWrboIGPT98mHfqFIFHAuD/2frYIpju9190EkyScs97hOWmXC
QTUnAkVKYtGxJDb1DeOhsvYOm1k11jrTCStE+1Zo9O9RrbqvsMx445EO62I6gAhQEs9MOpksA6WE
RcPK7JhS66wNMRv1tz+qFyPgqk2AiJtnOhQGtJZUbWN1hMJZo3goEmFWd/5oc0QgBgxDaFa6RjQn
twbpR2M3DCZuwP+D2jWi7ze7rsVlugyK/naLFSC1C9RSpkUH6/x7Aor27988pBSL9qhXvIAwAtYH
BowXi6e6+6+tZTIgbEn4tek+DFIbDiVp2gT0G69h4pbAy7gem7+viuWgMAc1esR+gg4ZhUAVE/Rq
ruSIGNsJrRYQq5uO//VYPwETuP0XBGzmoQZCJe58k/4OuShKq/uSD1Zhi7NwzRc9mFXAokJB9iPa
8G6RDLrJPwU9O/loDbvp0P5n6aT1wiK2zoKD8gJTkr9hP1Y4JNjBkFaxABwKREZBgMtqNqXFcGmb
B/2Q2hqkDGW6HjAUNPrlNYpOEEOrVhZRMDJcJAhcakfkVk046qznFwHYgcSZGMXQLrEM7l/+cLeG
Ax1+JSSN+VlOt23L61vU5u+fnoVWNkQKczteW60G7SGuNTQC55ng4KQhDQVXh9MGHS7PB4PYjloR
PmhRxbCFNk2tmtaf4bEBHAHs8+yMVfEKGoZGTUWGOx091kw5Frqcr19DoNIo7EcU4sPqjflT7RRD
E6c1QDlujXJLG5zSGlnSZvFfCvtBWoeTEOLAKq0CHDI9fBnMOThhdGYxlo0XKp2q4Hq7jDGOZWLl
fsVtNrAtZXhCO5e6dvXijpbNkc2xXUh1uCXLTHw0oALHR6zfo2b/vmS8ipy9NtYWOns2UrRPJvER
JpZNS/wJ2GWbIxbrMGpmlPmEXbG5+kLbLfSqCmmyTma9gLDq3IgMyY9OKyFSNZ4Ye3iEcq76YdYR
m5asS9cJ5nDPfzK2oMnxb94TVBWHfE/aPmhvm7yJqR40u3yPzLMZsKEAg+zyBuLkA5X+p8rrXiKL
ByjN7KidJ6D3cwq1ucvtuohO8qvDg1+M9Zv7C23SEfyh5Kj+xiY2ja1qRCTC5qEFYAVsD3bt1yfs
iMMd2hfscoK0tjq+uR0QCKH3lbQMLlc8/IJQp9PdyOxaO8Jw8OP87jzFMjZA0VAUXW8a5Tt2in7R
iva5pA4SbyeoPWqxYlLj3zxUI9RF4Gai+HOdkq76yA3xpxKZvX2jX5tNlhV0rZn/INp8JUHKXi0r
dpUJKRkKMEkSHGLeEl/Uj+7+cmSDF7H779ptfWPILwGv8ubOkcHvnXnon0J9f/2rdLB9disWJ6zE
xqfVYilTzVmKAgp7dUgQTWZTGE0E88773QwGyQzXNbHj7faoTszHwKObhdK35sSmFBIxM3BO+J2v
Om2/YY0XgrwAsHUV/5ha5q/iFiS3j2SdP4lSPIUQrT5ZcKZCuypV9xT37INUS96MrZIrpqCpW6RS
oSHw1hLilxDFpiaX+RJIgSVdxVSL92Q+aoN45PIMyNVlK1ZanJeS7CwVLXohSiWNH4DOQVUhj9BB
UBBH3hsMs3ED60RyXnm7b/8Qu0HpaSpyYqo9YSiyeJ1tlVXHNhfawzrWbn6olejP4ZgjVb3Pz+xR
RpGTOpGiEv7sMIv4oaj7XlCtExg9LiaiiJI/9TW0R6v1TrvW5DQbP/XaitmKKQUKN9isOMV4JwCb
L6d3wK9LBPSwHBWkKTFk1gH62IyCIxk7TWt7Q5f9ykN8f4r0bAxOsdnS35LH29TgvIFpsDgnZO1X
mgnFH8juZ0IYmgc830xxTo4eOGd0bi4cIj2qYuFZPnJpDnX+dT/gyqqSmepwkpe5gXqJMc6p1j3A
3Mx8f5Via7GGd9NXuhMazX8tnKprxHcc5yqEKfFL+MP6GzCXW4+utZNumhr6GN84UX8BsyFP9MFK
2igoCzQ9VGrSFi2ue2lMMn/voSxagRnZ5P2KWTZB/wbpb3Ue031xbo6RGjafuykEViFAgKwOG6jI
VlpPl+u/G4hvvUyskaFuWLxmNv7gJ4mX5TZn7jPiz1/vtlvzseymZ3Vchbb35eYbHVTvgMnMZPX9
B4WPpYC+VXsgGX8oWzlir5kaXb5hZ1lWrnNfJaOQkv/0UHS/LyxZEWEcnoY7K4BOFBrO5sF0kt2o
Y1PFRYlshm7G/fIhTo6mtEzaPBetQDOfx8v47ZfFXMixP0RT9jyK0zBXHIlQmzKhnTuKzA9H1vCn
J9w+pg8stMPqo3NJ99o8s4zHQNfaXfVZ9hO+eaTPY/fM++9GWo0N/IBxOvANwkFMdpiKDwlOkfWc
/g7hYGrKvlNUp/tt+nGKydJg6PcrrIhBhP/XJ2xwxwNP8f32VLSzEcCy746E1woxJn2dLnw4h/vg
Cc7Y85w7XqFvGOW0Q6V96EqdkH8vIAMRrrSXfVG9BtYCRkmPbnXyMkOGyaVoxrSS7bAFlKFqY0zd
CBMi0B25xvjsLPBredaRzzD9/7AqVxvCEeYa/pqhktcQOJwuyhbnKeVtfbB1RMqHmFTX/y7QWB5l
sOB1mBF+A47L3TMtl5hC4THQJWt1YOWSVh6bnqIIMF7TkCwe92ftItRJmXxqlpBb+KNQoJqT+GE7
kEHPOd5d59t/t8miSwhcDj+pav8DqX8P4L5DU10i58q7DjNc0uhP//ySxlSY2M195BfZSW75gbT7
zer5Mj05g53335F9gDYkZUGvK4PEIE8sZ6ac7hM23+zcVBvYd7VhNqbsHr0Eulumgngf3GqOZFsb
OvrF0EX2Y/NeT4L+ZKDm4D3QhD4t99425skJWjEwZV7CXG+m0bQWQdGr5Q0UaeRyCsPBAXA9eOlI
eBEpIRrXg6h3Km+Ime0KOR1wSI0xRz77ogjACD9CyI1ZwMdPcKKtC9vwQn4Aijd34LB+XRO3dm19
4wHBLq/EqM0TKFuMQdoUVKGQcbtkoOH0hmRc1yqLNHrYnz9I6QH0xIrviyAWJ7tx1O9CfDZFXmtG
Vd7I0QcAAoieQhuqleMCn4ycDwTPGMqHG+Ph9nXMaSf24ctTMrh7W9mMmmt2rOmB6v+7PB0D3IA1
HGv3WIe0U7KBUHQc4XZLLvH0m/2b0XFBGVAhr4gl15gCYIygarkjFOEDaykA86EcjVvhscsnlFjY
J+SEivVf8nru0qM88/DKOP5kvW9bSONJKiLgR05TyoI/QF1zvbF7loygj+5/wdTHrEbwn+Pz3N3a
D5BSx1EFqcKKUaCEqYhRnXVgWImqZucDKoET6xawhrZVDJL6KsQWhddOB5a7C9UQgyshOtjxFoGU
dlKMTHOAC7K+MqahZRj1bih8UUGvqouK4naN2IcpyHb3WWXXJzRHhASbIMAwBUi4VT35RbHHkDh8
HyOqp4VLQhcOwFpSsCV5cQsRgx93HP1wZH+m401dA6M/ZX/RdLZpDVtbaOqm//SBufx69qk5XvFA
7EL/afSVVixS8JWJc2T03lN9GtXXBS2zFy9OIAjE3FSKW97B/0Y6rRIbzka0XVH9CMmPYP6v6Z1k
XunRVtA+B6InkyTVCmSZs7mFrWZjMrPsnB7aSHFXX5F6SyhQ1D4bAZp0dmq6kJi/ey0BnB1MQa26
2BXln/7q6eF/RpfJC0RunszbQo2Sm9USkPb3BXG/jlm9SNVELKvWFXEOXVgaPfYMQoOpo6s/S0T+
1+OLhfVbpyw6bjj2PAMxrZm8l3AT0vYspm9awHvapQvX9pIKKm/VD6dgq1OAaY7DUGYpj4O6aLwZ
JQm7Xd+V7uNUCjaSdIWAAMP3BjyyXHP0SW8w1hCmlWkSQKgqoL2sZACeCcNcG3EarYvIEuSZm0Wq
8H4LWbFzEArmTCjx8OdBe86MbXAEcdpvhm0ndQ5jTlQ1NxoF3jLWA1AJYaml0mB6KW7ys4CVxvGF
tRN2/KzPuw/W+RlPJ86PzOy7l3jc077hMjHHy6O+lTi2Ke3/gWmH3AIMqBI/Zln8AcugeCV4YZpR
8L8OSf7heAIdy19/vfuyouA158qZIbY3gef51XEopDVY88fQV8pIDbtICkPMtIs5/itqXuItXpQx
QnlWDgBIg/2BnbeKlpgumd72JquHclUqAlTxH4rHRry7gSxm3gsMoNuSLWPOX6UimGKrPp+cDQaE
RIFNDW9bsFWePXMMHZ25Y59sCcikgmO9ChB1WoS/iS8M3Pxbtdfl3vE/9HThYn9hvgZjWbUAJHfm
dfzthveKUDvldNzkvgG2VVzhcz9KjRtjLhBQvu4RXB8snz2klu1zzPD/HBhtlP083qJGBqGisoWo
08dDIBZdG7cp0EDihJVG/2DLVJVpOz0Q6tJH0QHf0g4oAyFvZjEDLyxgLSngsTkKbfs9qwKs97us
8zC4urjMEmrZjSyHuZzGhrnj2qy4t4xeZaCBk+gYCBftUA4+JgzP+P/JXxU4HfxOGVBsjjau8I19
E2p9eKoH7ZRQRXeJb0J8/fnVcbb3ni9miiOmZo7nVuKsd6v8B9Gbx3NPy5fvCMDjKdp/4O6RYX2v
KEta1MlKtR6Ui0XJOgWGi5QV8T7xlBm5XepYDF3htP062w7Zr1ZErwAGaRMQsm3E0D1XaBU8dOoi
dNv+hBnPm8kcqIMqr0iTh9CDj/9eLHgDX4sM7ynQMvKP7PLk+bJWPLW4QOS83Z47McGuzWhPWe+B
qYz35jlCQKA+/XLwdZpQn0tpYfk3qgzN2/nKbRUC49twIUROEWEohJn9xjnZ/LLnuF1JLd1MoN8Y
HLF2AS6A1u4qQyrN2uW8m867hSBpEtg5erc7CboM153QwyT64Ag7ii3z2yekxd9T4I2XvD77eRPo
un5OxFPYPC4Cm2dRBbwWZDBM9s8JDxMWb4pK4Ue5ZsBZF3P94ttQfX5jERq4/5fbCmA74xMzZukK
RxJgpFYygWNKpuU4mvDhIEYsivWIIt6Kj8zoFy5uhaAHDD7UGF9xSQe3+KUexveqs4YjKqA0AUIJ
4lm+T/Cqav8PRKo3H4oo73DDqsJ/DBCr1sCINLfQZyTpPeFzMaoee31/gCw1EnfjN3KvyUAEHuXq
ko8lHIwI8ck8q659ACqXODd+kcLpA6vFHI2v1cVRhiQk075hxAP9EM7VqXGuaMghwuNvF/Nec4Cd
PfX0X7qgceneHhDS9fy2UihsAt32vKUudKLgzRJC0SWA0WmoCtXtBrDy7ORY9u6jOBWYtGu/7Rum
eQmkkBTd/SKdBBhu4vNWZ097QRMcLzzOrnastal2AuydSQGBgO0lCOGaEqaX2AROtvj1GRmLmmQX
IXhfI97nkvWaqtnXgPJsx5oNlg/1yziCmdU3DymhWnKv3fP/YsWXzEVQRUecXZkDdwzc8OXTxZQx
UNoZD9jBJ8/Dj7ISp7OmntNMkhYr8PLgn1FcbKlZTrjEqedYYLUN8x6wNHxxePkv1Y0Ma/Biu+zu
HTuuyd+Gh3cBpEIvI6PBxEDLuF+SLLIyrQeLtciY+QFWlgochNa8ar5jZP/uQaYinq6x/LBg9xrb
3PhrmVv/BiPZbEa9XO5Hr9PHqtQULZytj/W64MKz98/R3j0q7Ecq4nDEfT6ybZwk3j5kNYTP6bdF
dG9g7g94b1700Zxtwkdxg+UAqJaM5OAEm/ABgOmWKKzuwnI/KVnnFmXAG3DAfNdJ18H5e4+aFACK
ps5mY0X8HkU+wnWJDZhfjPTv+icmPW1k9kYwpCPo4pXbqsra5Hpjh7v/2FsF+s8p3xiJy8Kx4iAu
KCblCoNB7xMjUKyIWUYYl/GgtJTVienmq7w2nZdRvRLb2RX3Q0unlcJGYhrAwJqRGggFcE8zWcKN
98xwDn7ax4HHi+ao+o1od5/nGHCHH2QU8n8o0eTs8WaRZioRLbKk/xXFDNYQdZGXITgQPjlFbnW3
m2mIaGOKHhXEeublV+dNi1kNilHFg7u/m4Bdg1L4fonhgWOZ683MbZwNFM5qSyhvpfKJ4GXd3Vpf
4eVnXwC2DP5LSzf9bNvbJjI8V9aquMOn4lK51urip3ylHHk2i3f1PKgGHXjWOB4MLrpsmlzNp3qE
nA4JDG5/pSqsW4QOKx1VU0NQOWyaPieXrcnVt5npQxUb8B78j801xfc9NMO41tJa9rbghERytiCu
z7aQTsxVt8ULog5jauBvqAQ6f705a9FTa3BPtdXbkDO+9DWUwfE16Ka5h55rB27wxWltQxvL7drF
eH1E57FRxI4fhOR/uc2YYjs0/tXy4Oik08iO1GYjLTOnNcGMsBA2PSNmWWlA8x4yOQC315aPYroz
xhix5ixDdsDVe4+DTxPsPjpcuEc+J/KwHLWCc1PGOQrTqMXmcNZqfIc7q/heOrviVTpH5RWITeQL
5RCcpB5Nwb6crnJFlnJNT7/nfO1x9RE6g0kX2lllq5WQAG3rOksuVzPWLEweY3KopgxcWJol44pQ
e8i818K1/kAiTFFe7ZixbItGL0ZIoGijpCUOGPRCU4CghuBgpSMF4Yv9y/UNS+qTwQwQjEPyzg95
qyCW8SZyRmSN7YgJWU3QWOipBui9zvPBwnsTjcYkfiW+YgG58wWDS+82uogsHwELxAkP6i94UefS
PShTkT1EoYOMmWhQbIYHipiwK4Fl8TlcF3FPPDngZd181QcZukMJbRXin+AizYBcjb3kodIiHMXE
kChG/y3N2lSG7ASvZzFpACEPtL7800odDQJVBhCHIlxD8iy1ZQmgPd/nyTAmoyf3/RqIYy7lWjDC
9PA6to2yYsBmijC7lne/AdjDcpZA4jWzj7g9mloFwTJD87WEEwWC2jftL9+x2MonTqm/7z13TcKE
quoFdVOhY1DKRmmNQBMpUX0sp9j2BRHr41Zk0CjhJuH54fmmPbOPTNcWvb1q4a2KGLj4GKJqXB7X
RcF6piGUkkHfGwstxLqaV9B7OSwuw4jmC0ZNyaew/eZNEhD44ZTKV6shNsLbKEvdHC+czz15gx/Q
4U5eoQDdxikA/35H8FOHau2hoL+QwlPheE564YgpEyF2cURaVGRlOtvefIfO62bBPr7UFk311uTp
Y83E6DO+H9msmxCHDyOQdgCkR4yJf/8VhMQvUTxcrIPGAtkbrWlN4CoGWiR1XT/nTsAMYDKtnT3c
ikqL/YeE6/8ZgXqIuitw7wlJlxH2TB4YeHtFnvwI+F9oqc0fsQaqhjtpPfcQsyR1hfhqEOvx3CZ7
CYwxUY0q2K/YNzRvhZ3OdzIc68wC8lB9jpsZbczJkZjPW1qN/X/RoL8wmDUE5ckWnWzHo7+kOklr
2aG5LE+rd39IfVoNtwoelvLOBp6MlWxMp1plxglIh4CZ6Hcyjv7e8B8VMrE79wHZeHvhVMCMkhk5
ZGnp0+ZojyTC+zTnHbNYXjrDP2UF33zGlqJUE+GHLYXcf813ESrvxiztmc0CSaLglkvU8cNxNvlm
XUj41nSxosOkxVDyGzpRRcF7JwjdnTx+lhvPAZJ7jBIigk1fNSNMHhvuzCZxlruDwCVuOxpqqXTz
qrjHE+wabeu22y5qP0zZ1o0lnCW2uQig9sziFeVYsLFAXRE/JAZ0oDVD4aLnYnSjm6Cg9rQK9VQI
HLoi1YxnKs0GS5h6M2Xb3KNqwuutR4QXBR5oXJzwguevnsarmi3mSL8nJ9tW3lidAIaIt1KS8Eyc
1yV5vZHighvxb3vrIn4Ik/dOefPIcnVo8m6f9vLecngSNoumv7B+SN/cBV7AWgSRxh6LerAtqu1c
pLvkvVl0sNcb3NSakDwF/VCmqOT0husmM4AFtDuUA2QRe41ACitEMB4XG80xONL7HEbfauYqncMB
ScY/3ADsNqLYQD8pa/KJHyOMDGh30vPOCiqNG8+I0rzksUc8uNGHFzRDj8aHUBIAcnDqwS6+b/AH
Li+iLZhAxgJqYU9wgoTlIGgG+LkA0AD1kpYxiKPe8bspnqfK6jEr59aEJBciRq3/hSEfG5e7la3B
BCAZlm11SdikDzYJn4mW0wqpIgdRmzb9408WtKYfDaNNHm3eXagt6AR85oaVj0H1zf1msTW4dJe0
m+nl85Dh8q1gyiHn/Eeb53BWQtO31eLO5phi7mMWNzSOlxQbut6jic8B3tmHvFnCmJuvggP31s4f
/Q5/Ol0dfcJVkZXHNyzDmmTP9Fcd9D5/KfrDiCeQ1FX1HOWBgj9RkiA487z1wuEhZwAadLxh9na6
06ZEfb011qvl8HG7QPU+WSZCuMjCKvHGk87GllpCI82oRZLkQRwGwy/z6UU3EVLelv5lq1D66ttR
bbsvbb7D0v6jqNzdxaalRI6Os5eYCr0y5Fsyo7pNb18zUoAwKElewUd98C5M21HP+HD8WwcK+1cC
zfTb1/wZIN1jUHVErN1IlxZTYUYCDX25E3Xof597dj8Uzvt6F1uq5h+Osph9ofye07PkByrYPvdH
l1bWFIEFSsa+P+0niq7im2pI0YIfASsiFi+of9sZwjnwEzRVYwmgPavmkb/pGs8U9QSJbiqKuvUh
BcLFg+Qbs42BaPIp2PUqfvUzTSm79+2owpNx29SUqw6O4//eAnjz4B7ok0MtdWgFyTBkobIbhvJ2
X0mfjjebe6yaoKWB9g7+7Z5GbDTNp3bEVsU24Xp8BHEmoQiP6KNaWitnerG8f5wqbaF/gU6Ntqwn
lZRO0GG7kDqnyK6kT8qyDGYFr875Q+bkSxFPniKnNZTBNR8v+VvI6FmAowbBFXd2zHzvwFcBiW0E
UbKEADnnJ17XDKLAw+wGSJyJqN7WEPbIbOjIXvvwUDy3t2eXxFhDUNDnUfEG1iDSQqV4M9ZFWjam
BxjBsVC3RIZKDWhFGEaIqq0AdIPXgltpbX033B+OtduK8XX18yrNOWmoHZOYmdPd5RPF86tpLEAG
87mVhrADSNp2DksyHo4UwqkHnLfOBrp7j5XJODussfbQGSC6VhkIQnkcMRNnj+DpVJFrPVfXrgzZ
0XMTntw0KI7vHH3fsKiRcNaiGfa9Md8yYoh6l9V/Ys0Z4GB5+EO1MC1780ch32gGzAYSOGIwZuSY
uwVdJ9SyXeTpzmfLWlLyVnl4EiW5uTgALupg7u1JgXwb993r7nZqYdfX29HMydPUxT3XKmKtneky
V0dYLxUoCl6FxziyMAYdIUiX6lMlzYFVKRGKdOLLPxYJ8cb4Ae749ICK9XWDFx0ZPegQdp3CMrOo
AwVt7WgkO3xQJtgaLbG0MkjRU6d2j8KoQNtp2pKV9bvBARiOxB+aJd5rWCzwUfTxa7nMIsTMEr3b
V85RMuD8l/8YSifelpb26liA8SkCLFDA80D5LKB5SxvmKsY0011+6M66kb/kiHyJhnCk2PEbWtLt
eCDrjwzAr1slYPh/QV7bE6YhSrm23QruZQRTwO5TDEw14cHfG3FTOQu/XTpGPkwfBYD/okIXCokZ
BVbInsidV83lZyA7h3Gv7Q+MS1AyI3MPp1fheevyiyzHD6hnziDC8azCOTxwSoGKV+g77knne3rb
IBifNipwulN4iorQhBWv8iFFX5Yun5FoKljwLh33kImg+CeyKkewpeO/KwftST/+sbp0EqRwj+JA
spqvZMSjYWF/9L6rMr44pIk4KFFARjT7+v2bp98JVqFlrJxzDt7YPeaA/eLo9aN2WkjgT60PJWyD
f2Q+QNMlxArT3RKXg1SgKb9BYcaftchQ4PKZNUE32lvV38jJpVKzDU5MfNRS8gHc1qPqIxDEBOBM
Sk2q5RmBT01nwMACjwL0e1ahHEt70lmKz4FVlAfpW+8FAE+6b7DsiVNhyDxIa8ZWB4KRcY/WMDkJ
hv0oXq/FsdEQyFI/cZRWGBVxGgDlmWotwXSbMnQCiR9YYFxflZO4qjKDgIT3sRBcyjqImyRMcUqg
qPGUz0dP2yAlvj5G+D5qvWlWKV3EeYx+QGTnOIbcc2+wMAftJ4yDaf3TrhU7Ag3b7In0y8Fa1oqd
fqZkIXm7KFG8xOsi+pJZbGz+VJHX3Z+HcZ5uEAeC9lYatqrcJqXaS8GXMqEnUZPYhB4gXxnqetcq
m4BCsNyhEl24RtKAy9FJtad8VGOCRPyl51wCAcb/YbXOmEuD1SMS/g4p3zgOyp+bDQ2ilCB4FXcQ
HPyztC/GufreCgBB1i8Ii0u+6yuFCWETq44yZ6AfhcnhaBOBD83o7dOVcUdFrvBkmhchslqauLgC
7eENrzYx2aXixctCbh1tAPk7WGQevvLPjiXTGsbSBGxYeT9qW9n6ZDYenCU70S+/v94E6vI8FJKU
/hcQqOyNEEiqDVavz8arIOI6x5sF84OhXaaKZ7ePxDOy/KCxLVxfMHamUonNkCRUNtJfusB3sYbx
5fOngtn4dbD/Ku+iMmEkA9co/UUc0LV4wJcoJsyhS/s/h3rS/etAUDbpbP0w9HyXskOAsMvtQ3/J
3wdHenT7jTUeImquRbkqUFgfiHJ1vmjl9GBBQHQI8HZnityW4GAZW/jAtn843WPaituOwfPGop8A
Zi3oeLpm/NmE2IvPGTIy/5aqt0Hqz6YTef8qX0K2Sh1FUo68GvewG3Rny79eIx5EOcpqTDp+37KK
bCkIf0U1RhKssJR+VYyZG4Q2AKcnho6M61EWxWgU3PHPhsu173iYxUR0H9rgMPsWEayRLuOgV1Na
/bMAMd0QUj/1GhhYNCx6CvnO/Z//JKLwJ6lY6O2jPNgFEuj0qdqFxUZ5eNGfucjI3+5wztrbjerm
8r1JVTxAscTfMVYIxXPWDu1UG3AvjNZS3KQL4+nHQUFx69BruIJY5buIwWuGldxx1SYyODiryegc
utAwHiLT1b7CfBSmj3MMrHy+W5DZJK4hzVGfVCieNUJMMpw8LrRfMvoKlI8GxMwGo3NoVKhdwyfn
dpXUIsCySRCnbKk6qWmsf55ewF9AhIu8jX74aOFOQmOeE0ob3Nzzlxudx9XZ0nxFXir/PuslF4wM
hXU8nwyZckRNBQOHR8KEf0EanGCOrx34wB4a+uY4t+nr2tMtt28FcP6lBHW/zNfELP8w7C/9RZdm
MEC+VX1X80QkJ56pt2ZVZKX0LXeDie8jMwLgpxO88CenDNuASp4GzyYYeD0H1slG+4gA6n56LnJh
TDxuGi2aQTemOsSnFVUL10JH4SQLqy2DHkjEKDr7vnUFo8tO76PFJYnuVo0eh79uTeWdoMrSS6AZ
HGz/H/hdizPSomDfPB83V1OhwBMYfeePMOGxgTwsiOUPUn2ZBVVotpxfSXvyjiKy9eOcdgfBNFTM
xBedf/tCbq9veSPxXvlKoealDnvhMbF4YwuclcEaEJ32vbh6FsQ4nSfJrX20JBrKA6DCy2shtTNB
yocYwiP+YHmJa3VYVPkzrocpJQCi/B1uQAGBnUhutWyHuPZnfVpwtaOWU0bFFn3nkO28+Rwc9+CE
qev9Wfu3bOkPLLMhHbLzyM0yXD5CY/+EyrpPH1aC7waFEzLfTwgxDv8acgKx1+vN1PSTbEh2xze1
kAi7C4PCAu7RJDB5IZlqULvt070b5Rn7PXmmGKuj9cud2HWcrS984J4pOXJ8Y0RuR3O00FlykuyY
vV0HvqAlElj1k/p8pOUTLGaXpRmpmZ2mUOljPjwcr7rsSGoaZ/4SJ795K0jX81vPbC0zCPduuiqM
RHZPN+qHkPPTCN3gmh45NsLdXNsScjxWxDBks78rkbNEqc0qRRR/BQz/zV1GAKjaZRwW9IPPPM+F
+jkbjAnU0hDii3/1uf6jEDg6F9Q8iu8qcZCzZf/Foklt78ngnFVses4/B929t3My51+htrUZ7bz1
XwTk/rR9E+Ysr2FIJQCED9pPWEzMYh3AhiWglp+/rwJERxStZbR3R6c9UnzBzqPZDqRH8zHo7Se3
DLCNqHfz3so7h7vVM8Vj3xpGPY8PHvr28tZT2xvRVPz9vmS2Adc0tMYcJ6PDCpcYnl8DlRbJsj03
iYu2UkLJpckGZA5RqkwJ96K+s19kG3KsjtCPXi+5s0Q9iuQwrCcbPaiRBBP68hK0N3vMTKsD7qdd
EX/k7bW50SwJfE3U8LUIgDDArLbVcpLu1+GkERQwd28BDQotzEd18fy5SFTCLExnk+H7+lwM5wIQ
zk+KzOVBOtSada/UO5FIayEpre3iZZpQ6gUOH7KPLoj7g1rrnPNVPx6TIjYZ9fUFP0q9oFIiO9mX
aG+uqnuU7UfjljrwwrQzOzHyLxk1otsQHIhXuQhi76Yhzs1oCZ6ykKILQ3kF8ANkUQ7d5srh73XE
TGN47hwMh5WaimXaCrXhf3GLDtKgXJWwax0gv3sacezgd9Ug70uzvPH8m+xht2S06lXVMEaoV8Rr
gsrZFekRVXTtWXzMd4W3NN7YHJiO81PfZRDlU5kubxsLxrm+rRqrTP8SheKCWGwMRyOaIl3tyKVP
AxgUFxhQtrk5/lsYwEpk5jH+SDq45wq7rpJYL5fiHin3qLPzR9d+1pInq9fXWCpDM1lysfzG6kFw
AjrzlUFADIfX7c4m9vDYMy0x2WZhiZ61rcx9xQj3BkbDmp0WdXMSJ6psU0dYahQHa7Dh0xtRTEdo
8zl5M+vYAaocp4Xi2316rwKl3plFvWr3AqDlVm1nHLxI6IDD2QdONmgj+RYGodnw/9oDODY7KCO8
z6s3uvk2C2m23BCTS8LSY+/HxHO4hMz244rEe9NKxYsNJQ69eKh9Rr59i9mKTH86uFodJtEFXZxI
HrGM06eT0aVJw6QCT0tVZp9FaC48X0XHwGY501b6uMB8V1nkI1JShzhXxoIO1oyNauhNuiI2ShC3
zK0b+Ays4epx5Y15ALtMIluKvBhxKyXl7EjP0zgjMxt3NXG2oAXafctJUk8AgvDwYC9IqJS7zQNz
p1usSmSXmz7/1kx7zjbS5N8+7hpWtqIumWNj8pjkS+7NTRw3AiEXFA8PiWMTbgaogAJtwKmhhoE+
pYmapBQBhHoEXNDNtNQyU50Qody0+V+RW1wnv7kX9KL7E3Q7mAbaV/5AijB+EiperyLbCVue0Vtw
bZscS6itguFI9raS4Rb6EG+/MAiEnbwoaFgWFgb6xQlNt2VtDTPm5Zbkcm6mxQLHrPk3Y5Pb6EcX
N9XB6X1dgAMdkscv+d/zHqSMNsgEdHOxjo8GlFlIzuH84vXpl/XkJ4/fRWtllrUgQbUy00mlr7c6
fQyFrEHc74NXlVfLXo9ZDX8TxCVXB15bBHgrQKHh2/ZgkIWyY9rH65B9DCC7Xmt/E92CMXA31Is2
zWik+AatZ3rbr2H06ovpSnzyW6LzaLUzTzoz3oFrq41B7tIihS8sCbCToNth0T00UQWQORXJz2IV
76VcU4Kc3dtDOc4j3XWrS54Shwr2ZI1LTy7gXUWISFhWuzfhyQ8AOZQLAI300KUI5nDlPd97r8wa
EuI9u/y2r+se9FGiUaWBINv9e5BjFZ9ZpHsuDmbSWSTUqlNGGFtpZBKXRXZBWuzWga3EAxHdZzew
zKyD6jwFPohNI7Zqz2+IhQOpggzCRgHOjaloQTKTIsT1yIlzAHE0lsrtRzh18fJsdlYrjmDCb0wN
L1VznKhvXeWWX4ch259I8ksAoKk3H5YRg1SW4rV5dzjV1JYt4Ek8o7PXHOmMaxVzpLObHUwJfDOH
VlA/SfUo6W3qVAqynTAQi7tb+IgUjAxAPOWtv8vKk3+8DkO+v38p0snX93EjP57/6yzhhsyQC7HF
8nkyQ2jVdBQsXN/Z+O1Cw2+TUuwEn7eRZ9XA/WiG+2aKkqFMr62VY8VaaRlQ42vbWm1Cq9+emVDY
nsJNtDjDg3ZdQTer+MLiZhNEwnnxIC5FRjhvAtRmvde9JCwniX4RwyDilRkHCrzLH9gH50a1iZvX
07qxVBfGX2z3P8+l3OR0fQSj1cue6nSWSxKLUImmPeyk1K9vdTDx5BteDZj0Q0mK7jHS+GFj/ffL
M4dPLaTuREXuAAl9DY09BVCZDFNqxqtkOBYKfRIlY86wlKfv7B2L+y1AYmoEU5W5RzoJWRVCzlur
4SHFdd7+ftp1HNad+oMOJ1h6adpbO11G7NnH8fs7mbMZEW0Avi8qCPTr1usbl3qHMBoUqbQIsIiO
2mw3nxQuvwP4GTLo9hgaclQk4gaAbIoG4A05mlcqG4S59A2M+uxS4bGrWlPEA4egbJ8LPGZyqYJ1
V7hI3T82idRm6YQt1eVBp3eZpBsfDD94Lqn82nneTtlArznfMWKyDfHcSu/Tx+zQ81cFD3i/vKQQ
E5SEj2VHRqcG5NmfcrCAb11KPIThCJMGDuUL1HfjaAjYlkWgOI3VsHoHqvvR3EWi7YwEmSwDnx4n
3RqaBkO1ocD94Tqa8v3pLlHMiiSjJNA9YYnt9K6Unprn1VBQxKosHjCzIXtQ/uBqZynI3PWuUSx8
8lEbYOHFkrM55gNGBsBZg3gM/+P3pXMkF9nODiJcJhoiuAJYX++ZUnuR/bMG1Fsq9J9ugdH8cLKI
wteXlrtgev188ZZNIjkBPIku7jhCtAxvVqJ5Xq6g+TWe0fqUD9NguDr/plpPkGhDPFttcZRl2pT0
YuUI1u7mvLBzhNs/2srO+whQ9sVFhd0TcGsBrPNFJsPV+gdDRfAUOnIdidqGwPAxvQyrchltGuwp
3DOBg3u4xMOmBRZW0B6W+fEA2ahBJgeWs2BiQYS1r7qKXErsNr7Iys7r8Z2Zr1vjqd51uy1Xj2BO
R2yZIQZtOo+0a0wAjc2oZN6Anfm8WDM5DGyWmw2Byvup2s41y5FwDaAYQCOv5MglP0KGa2pZwyGP
sit4ZD2DqQmE1qWtlAAfHDMnc/GUOF8RvYtaS85qqB9fTzyYqV6xpMdtx+kyhQ0IcUpH7nvRx+nb
Pj59wkkgcMRGF0511vV3N6ILcMal/Q567hDsIretnJ2FwqQuoHN/RQfZxK32CKircXuH7JSRC0/z
sIVvOM9qFKt/9KpC25c5ypCI/lUi3jRTmw41Bu6xtUP77FK81KeyfwB/n6kKmi2cjI6vLHqcoa4O
4A9qckT1pWjxmGiOOrrZ7/L08iDkYQ9kwaA1qgAfgKt5LgUi0VBofHldlaM/VcOFdkOjI/7GfPBL
61VJq5kMfeipNwUdtLEeIR7DrilGP9aNYcceeRwRpZMZxEzvlrBoGiRgbzzLb4tJzjw8JhkJsrqU
fDt0bWf2/mT3YcyRYAHFXaqKHxdqDjecQ+2D1Nh+q7VZh21RdB6AberxKfSU+QaelpqKoW2P1Z1f
+wSex5KmX0aTRY80zscAie249AeesJqnZPA6MpZmwqI69QD4j70+32NAmsL49VuHsZFQL0hULNRN
JhPdnQbH1kUc8f+Zl5B3+U2YgwO4Aeaugvklj3Bd9miLL1Pe/frUerCRKGD6KxL+QkpzrQIXFPmK
NQayui9n/VDbmtzQgcuj/KJoQh8Vn0CG+avEHLP8cCvI4tDiV9e1IPzitphTUYhQ4YyZmPxAPzGS
1wU2rY/GGA78ngD05sMYQissLBhy2RlUREDTALuZgNxcYGWrQ9PqEGS3ODoy1WyIkCGviGz8r1lI
97m1JvD1Q7THXfE96Cq/WdC11QPLJ4Kolr6pqPT2l/dnIrmPWBjYDrbDskdnw/W41Kte0oH/wg07
9mxfKGcz8ibpGVf+UgrhxaqUNV5x1Rb3+OfuY3LJ0+PpJSP98koNe9WJNfU1LlGrPe+7sep/62Vb
qqoQj0wsgLt7UkHqXqVr8M1tgDwchfBnm2+ZSyTHzdIgWmV309blQ8y1R43sg1Zrbz8g4W/Ul+/7
AVKm42iZemvoebs0XWmeMR8SIwQadWnWW9F4XifooU+LkUnyXIQpoHFYDSs0EOkrMrEGr/+aMj3i
yhAGqKq45unMz52THvc92tdbE1M6ED/O7SYQJcPX6I33CL+Hy4qB3NhkUtRQKDk4QJFvwF6j43LI
finUkYV1gBqKq/3VAKMsIvesBENQApI1bhY+vvwejqnCN24+uYSeRZk0ViM+1AUtvnABBOJzkyc9
FpOBisRnH5JyyBGyFTUoMwSAoWzCUoieWK75ENGwYMFv3pVRQoPVMN6Bl6Dmqm9Xz/mLRBTKZkxx
vefkXolnhE9VtnHJpWAdPIYUcNKhBtZmmAW4YfSEaNoZJD1NB/7/6IwIb64Ofqj8QlrPAecyRwzj
CNf4TsweVg2U4ggE0X3DmM3TXVuII9xStGO8CFxeYzIQ2FD3eYDcumz0NlViolxFBkrEeYFlh5GO
jI0smrvPC/cmLNhhuebY8D3NBdnpFfznWl42HWsDWeU12DnLKeMM5jpPNmQIi4bvd8Zos2To0MIM
nvPOlyan7CSUrN6OW2afodLCJqmsIZr5Je9sRCYoHUZFqwMPHU9ePAx6VcNzNDQEXl6HYlOcPHz0
3jwUG283S+T+lbAcMMJLK4hbs8lQU+1DakC2pTGCx9wasxXGR1rVsxLBCR0qAGjYpDvBrQfwGngK
H/P2Z3ZwP2FttGf6Vvu6+wlX+q8px9slJ0Q7sJ8EOjgRvEtwuZ77Gasyrdn3u0phHZWolCkh5BRg
bp4dq98ERP4ia6ZNPblvqSRXGZaJpYCB3uk+jhSpkryuO1F7S24L4LeSX61onHqKwcNJxbsRPWuZ
9WLCzKdwmf73QZNknnOKqcNrK2Pc4wSiMcpkBJqdoxGHWesE7YEtPJI73AvJvct/iTTnCc81rnGi
+UNzXAPjk9N/4OjtFdjIy/WE0IftLU+EJ4ZhnEvx8NXHN/WRfKWknSd3qfXI41gVok1GdNQGlp76
Kk2B4TRNBM6ikrjvVDokUvBur7ZzSzJ6YPzlpfDHWKFnKbduHIHkFQinuy6gwSNEa3aE5rzGRYsh
7ozGKHpbP8MbDpyKOrHsf2pNsnhhJvAZ5GNqTIIDti1IjlOgBKoRkS3Pfe+l2t1lbWU1z0JrwPhu
WEOkEMAy1sBAORN3GCtZCBlTnkdoEWVnfbW6rrTW3WYmWxBkeMrxXp3AJHsCSVjci/DrgADt0yit
QEQ9a4y0e1J9QXq7zBe88LovsUohEZ1iJ5vZPSAnPieeN829b0tBEoK/bCtwH2JGebSaJL9ZiDOE
T24lqzLoBs/9ACAJEajlMfF5TQGqIviySm3zb8YBk1KQtiG+tkVyy/59RPMQ5509cTI++QjY03tU
Dj7a1rhuYhGTNJyXBsDDxazstRbtXzrggQAD5PqWvu3skxcNtbPogw1Cnt/I4562xlY6iFXpZu5a
JcwdzVcblDRqmXenxNTp0km+Hwx/fVoeCPxaJudIg0Kv2CqecLpfK+HZ+emIqAQvIDbxIrfh3zZO
ZTAnwLlPMJrcT6TvixoXqXHY8YKi6qxK/rdfZPYHH4jPhY1phXi+i1xrx9pHEIR3yFFZbxcclw/K
G43/ZFcCDG4Iu9xIQk9rOmN8fWCMK/aRT6M0R9BHc/t4u56M0Pcqu9ubS5A217dbUh4ZNRwfL0IE
oIBOMnAylkiMgs/2/mQaAvBZy9fUbWtZgoR9ZisV/+q37uqGQ05ON1SDh6nLP24qqBz7CN2bfrn2
TWNyoMp8u0j5j9dX/sxzrBn50X3f+0Q7p8JpFS17e9r5sTiQaJ9Z17oYxTNJZZ56j+Nsr6MiIERi
W5clOXqgeaQRS7e3U9UWiPxEAXjVGM3VEg+yLmSEE83h60ke4NnvOE6s0tdtWqk44X22+1Fc7PYp
pDUWSkKQ28EiKaUwGC55Xpz+k9V85TjG88Lp6jtrdZ4AFEanUkpn6KkKMSYu0Ch3vFZLCOpjrY6o
cw+vW0iuAmFuDRtLDtF0mBvREpmJ9kTXTTQFlKm/SgtLxZvxBdpTOCpIDRfzagXGzM0JX/9H+B+2
drW3Ee4q0L57HFeQ6IgeNamMG3lNmxxDyvhSDPLqyk4C+5YyeDf27IJjFwn56ddpGpBsGrxyXN+S
vcM8ReaM3MyUQcvw7DeO+/tiIOV3X34xgq+j6hgRUPIK1kueJO3FMxVztnHZHMrdZNxx9L2ZpBNQ
szUGxlwe2fCLUxz8qNTTFe7i8sgxSshNv2v4GkYL3EpaqTLStIm0taupra2VlzFCTQkWagr7kj6O
6MhN7h2dkwj71WffF8V1s2EvUtEzHS6JVUgg0eg0uijSMlu2l1oM5iC88gE8IucTM7XssVed+3wy
06k/UvbSlCZG+6ywpUVDAIauSlRQUr3GlrZgAmKWeKPnhdWBMu//bu8lwiqzTWqfV6pkuqR8RzBh
DiVyjJslbTg/+5BjJD295jxAY/2S7Rnb1l2B6p8QvWAudcGsUvJ7Js+xH51b8Hn9+o2Vtjko7naM
RB8P3JeOScDaP6knCuAFrJGQHyLkMQPmFe9IwrjUhbW5hzL51uhPIvN/y038FLRPCsThWvemzsjV
eNYp4PYoAZdZmnK0m/qD11GkXqJJgvHKX2FAtPNg6wT5Y0v/bScxsdKbMOzMsZj/gt1JRut/hWg4
TEJcDlt/6QJZ1L5Ohn+BdLVin5N22y0CRhYpEdwwbpKvixTfKx0j9FVgi/CNK4vVI69OR8CBsoHS
Sbv+02v5V3guUf+/LwxCacWFXTiPeSQnEi/2vkPNdG18zU+m7BNyCmVciHnEIYHNsgy5F5YUHDoD
D6huYmjYAvMap2McvQMEq+wg1kJl0qYh52DuKKSgsJpvxrt7Um7gnIjMDL2a7D8ZMoq4hoZsCOHg
uAymKV+ty1YujcbKl89xrp85JSdUA/jvoA0mqAi7YchW/m4tnLGapCfaMUf31wCya8fKvk1o1Nwh
yhtguyo6MgHE3NZDs5LOiMnMv8f7N9NWB3hEuXH67VnDAfeCxibQ98TePiUCJoL0T5IAx4pJIIOc
TJSsCAIRrYK2XyZALYxnAT119t9e6l9+4fNY0d0q2NgbELxn82MKaFSPXZpCE4oDCNzbvVhsoQNl
Io2MrBvnkHspstvAA2HHjGlQzLebDN4z8trlG9hkn/tHiaVf5sBDE6bohpTt/mgscETSk9pC2KtW
zLoeK8zQbOLQwsHSKBeh0hK4z8cGYSVhd4JUlhzJF2clNMGigsT2Ja9OVnYKJA9oIxi6StE9BRD+
UTL3Aqe4tG4sdcuPFqBO2ef4aNy4KSHo1TNpTMsi/evdYX9uUe5JiFIbxfS9Y6DpX7GPRegptW7U
shxPhjXQZAnL3vqscPE6IqJbdOsNb75m+ErjTsAUp5RIbNUTVZvNWtM2L/89Sybz7s9HMFTDHN7I
pXcQpJpCb78Flz2vLhCY9bT060mmnQ4Ukip9I3jb3MnArsmVYa2h6knpi4AQBC9/bWUToLOy+7tW
Fniqt88QiqJBbTsOsylYuBXG0vIrr1krE9siKpdiUMnCeJwSBohKPCU78qSy6rbR61VsvHMHU4sO
YUKTku17MG0yNDbnwycRw5oC0yY0V3km3aZX4nN2nwlcfxgDNNU3JhNAqctRl/DFkQFBvTQmeKmM
iL/5pUGBB7U4BVDU73XPUYTZk35oCvO7QaAQTl9lcPdJxC11iqeVo/2zX9pd0qUhifu1AKHWzyP5
RXzhAKNZOOA/tyrjux0yIMRWFH4m1TXae3pTtkRRZShSN1ayRhU2G/tjUTIyiI4oi6QB4wRy+87O
URsPRGAv7iJovVTFacl9rJ+Nbo9adS0cb/Q+djg2sXaqknLvrR0Kc1DfUlnb8J/xzaSC6F7qsQEA
WapVDqZmbLuhIE+30pZVlUu9flvN9Kg2ALiJRV8EFkPjlU1hGyBrZZ3icf1bolhmUk7IMqTfkyiH
Pg67gxf62y5xOALdINYM0koeWUMT4nTwsplN4tkkpyWp7OztEi6rLj4Cj9d0yRdZmFNEz7QcKOaY
dd2w1XWgqGyu4mSLEC5JcowQXt5g2YMMhAF7gx3nFN/l4pyEZ0VaeMdmn6zURM98q4HtiRWZRLQN
CjKL/dyy8K0yGg5PkUtXqyik/zzOcHP7sWFQRb4mgvsDKZ74BwLP3ntFsDx9ZBOc17pJ64BO5Rgb
AzD2Mw41te+5oE2FWNSGecPQEhWDybKZ5q6UMgy916nwmkL50jhi6QGEVrrDEuBDp6AP1HXSE0u7
dvGWOlx+OGzlRAIy3u54fEEZoq3y/Aeo4KknKqJknaulMUHmZKEzkXcmWKbyFr6DHusgAMGijm4P
iYC+Tqoo2GhWFf5dob+CHZlbJBAXiyCmCD6BZ6mBirnuumPiB4Qs1OdaGWF4eOgKcM1sPAOMkz/o
ABjFcXHSQTiTFNcgfOEzsdrf3xz/6wz/MAspHnrm9Y1ZPxyzH277Wtaxx5UUA+KDA/JMf6ieyXso
CId1h33UV8o3+dg91JF7ZV7uXzZX1UoLlCU0PpoSDKNqUkJYmJC+FcoQ7Gnb2jqUL6XrZbYFCmIB
Cw/a1wWI/3IpoPqWbP4CUbA2K3BYyFQP3l5RW3hj6+oYt9z9ijWnbFemkAEi8HNHQ/lXC3UVexyv
YxfguDpz2DGcWouLr5Pa5h+kJN1Lo9I+oHuJe6+DS2PtGgUraKmLyf81DroiF0RbJuHSUutzUth2
Rj4W5u7fj8FqAndyJYYkbYd7lII6j8UEIVx81v3xKB+zjXIOSqMbc65CNkTYIgsMSi8CG+RcriG6
0+WXOCLe9Y+xCXFYDO3H0ad06j3osV7KG+TtG6IT35amK9hv8xBFwiPKD6SrSiJY2uYVgAzYfiv5
rmWPVgBpz3MkrSUDArbNo180nR8cWocl6/xVN2MkWlvv2/84qUwEdsTGLmLWXNWOdpKryBpCnGpg
HKPRKTEnTv+iRrcHwXbZO+bs/koLRlegQRL6CiH/9bPSNLWoquy5b6tYlFbw8QyAPEECKRzg6oAe
u5ToVxbNhN+hObCa1VeZYAtXR8SRz9cypMEig6BhHO7JaBd/PZFQIgvqYwYPOF0pPgN6IO6XBwYI
ccXq5NmjGKydEv+ZpmKmHcsWeJq3X+PlZ8P5TEnBrHrQX4T12UfG5NgC2+f+yiUGeAMpETTX0QWR
3DjIcGFtkH98m3/g/6s9XzQ56yeBWgdGlyWTUiLcQfgkn7miBPqwgfAaWVTG6FWKIbcVQbfPvXqa
cytcuYouJKb+E7CysjQhto9VGJ+vtsPIy+E4AW5kZ6ZiuQ9CtXdFY2b5W9WWXNsmYdq4pQb9fJhl
RZD0kghGH6YRGbzJdCFmlYTiuAOmLqdHXm4wFht6EHw0QKrM67gVkR4+zXB067s8HAQLQntdDKrs
pki7g28dowwSfoTY+CaNOtNDTjLgkRtNXGx8RDKq71XknZa+9iRIT0tzP9ZVDVP4oqm2m/Wl68th
jQZ1aQVA4sOg0shsFDpK9M54Wbrsg8r0Bpj83sFGZTcby2QCx6IRa6iJzOQAiOB+oX9KI4+Wdf1m
JZa40FxvXpVim48fGNfvcVHRGVXpLHLQwNdf8FKfi6SCfIU2kdFwTKLJNkqo5T60P1obENCVO9/L
40trOtD8+n2wflt6DkYTC5LpxxWgzh7cygr93IQrLjAHgBGVJcMvJsUjwZxrZKbqQlFdjdLMOev/
FGhNDaB149js+optHsj3DbGwfQLLBjcnSk5vprXPIRk0CHLFG+uwqtMQnzoCqsyBQsWIkTk9OcBq
CZ8U/8I8FMYyo84h3ogt7whi1+MlTeJ/wwGWs8lSPlOAY9MMCgKCZFKTj7l62WhOwuWW2vsbo5DJ
9kK64r9HotQ5Pvmmqj7MYWByXVrnp0HNU41L5RTYhBrbvq5rauZO+6myKvsrED/56w0fJ2jcTaAq
jnToTHtja6pCh2B6idO5Ql2YhvUttUlxs2Ult5QiftIRqnlmLTPjYTgFdlOFPOU7MpR7BujcU6Ds
HpFqN1bcAeBkrtT8rcOLCJ+YM+F3LX17dEH3kZCjfl/JheEBvBc+Q1UpjD7OE4yoEbReRpNIXc3s
3cf2a747msuOjvl+IEYFHR1R7nd6khsuG7bHVEX+dy+DBOi7n68FcpST+TUCvfMKto1cxwhLjHtX
l14+pEgSNd8yTAbXo3t/lVF23rplNOmc/lsQQt56l6TtH/fBX322uDx4MXFwcQunHroV2jxo5kIi
SAFAjMlf/MeumHTyIhfmHAudvv/gFrmBW5nSAXl+mBuyLRqq2t8vy6U5lFgbBbDcBeURQ/FYX7gD
NVAKMbRiMKlgX5BlbCoRqYpmAttuSL2XE86eR8NHHT8qi5eJyGYrDA0FlTdRbd5dKsqyOqD35zpA
f1dcnxg+JapLCQ0FFuykL9MZXnbWgKKW5g70t1rD+oZ+7oTaRkRAwIe/mGTtO9WMde5dmDglwp4j
NI4+08WNto5z5XafnRE4idyJBm4dFShLZ0Th9NmRzzJBl4QHBe6aPLGHL4M3LT8s8hQ7jr+B2TBN
ad/rJe/F/PFsksU5BbWUY/+cxJ25OfC66PtAIrsmq18JFLxSbwtF983Pv5E1xb7P7o7U0rXQGOf/
YgDBV+AqV05yxbMdfSulgxUv3YRbV1+240HFIv/3gQHzAllwigJqOoK7cbnP2VSvPSpP00NLP70W
8iU1Q1lvX4voUI+OzvGtNLiaIAUrFlh9eElkl0AbHwA8Rt1ExA89UDUd0MeBrolu4lVuUdf6GA2B
zbnN3LDw0yv0HpHKskrGCThjQ+Xcu+E4TK4OvQBr+ULfxOMQ3a9TJ2tAxBE0/LueT1++ubTXdB83
iV4GmQyBnqOJD9nunZjgKIuh4/bMZgZ30LY65yUWWDy3qP6LhTGgnUFvQGf7arzCJCwFA0jftgxE
VSsFlW5qPj6cR3G54dc7mIu+upWEQ3Tn3o3ToFVtAUtbWDJ1Sy2npo8ca6JDvVgijFFcTtgQxUaM
jYdJKyIwTERl3kH7ocByizu17Vz1JrHfUsbkjFlz7WozOmMZCfjhBCg3+qimlPQ0hjmlxRmMBg5c
tWVcegdCfazx+S6n+JeYFTbW7osHzjgmhFElt/pPweKUOzHMvVdSkgQthHu4ayBMtPNZC2J54uFh
wH4+8Aj+X8xIovZrWHaXw/uoRwNmenBMFQl8X4mOYpPhkj+CMgBHWwxjNSQcrGlTJ/BvmdwG2wAm
/uQrDzcg8ZkvkGCwbONtRbEmnK4ph+c0Wry2rxd1dxvOZen0IyBqULWGyoz9Nzm778uTygtFs/IX
y2FjL+TzCBop0zB0/upqAQ+lu2iIfGGJs/DMwhV9+KTmyVKtxwbkUdc+Vt/csT+AXkk0PW2GzcyQ
CRV6Kir5LZVQ9aZru/qsxykUaXPsQljBVwCvIv+kqaJDew0xnMQAOo5mKePuVj25klwUQgjHbaDT
oq+isR7XkDhkhhvxQGSbnCogbineoRfhh2Jo94r3PluWk4bGOHvnyxwqJ7yB2KDccdpOeIBK9eTr
cq7yzJ32PS7e2/t07XlQM+fhxkZoUHGrGKPYecZ1U6OMypOrXYBwSNRbSTsJnE3ZDgxikPXFZNWv
YpSHJjs1rQ0hwCB98RWMIJtv+IN8SPwv5ifbzYrjFYc8xQpZGi+VnNrixk7nlNqwe3CjenZky+0r
2rRtxkg7XUhi9I8NXx2VpJ/R8I79q7m3G2mYkqWhP77LK5zYaukg+Y10g/5f7moeDISs+/pjO2Jw
71usojqhsJt4ddHE8hUvI8MLNAnVTOJjkpHWYMBYrB2ph8aGfSIabJ3kpKMR2NJBVfXXZuOarmg4
vuN0OWf+64wQTruHm5GUGRoxWU61mosiv3xmg23uvbE6N+if+fli2HtNB7pR3iMU+Ld5Eouj3joK
n/WzcCy9Xpxd00J8MUT2jKXwW0M1CbEbg2AibCDfemqHoFAo2VDOUNQ8X2Xdm7PjsqpLGQedva0M
2F+RlCDpEmxDbyg7IeQAbS3OwkwiiPT4GHqsFuljGWNJrqADlcQZjd3FgAAHdMv9PgQeF/WT6XWO
j98PeaHjNkq7DeIpmMh0sThjW5aVf5IqypNNTwiuHqh95QDKPbW8aTwPEIgJt4162KPfHB0pty07
5kcoCWJhB/LIhnswVY/HAsDgc+9W6tbnAOUU2qwA1/voCnBtYLrpSHi9xLTVnTvFjY6Ljy2hMOIJ
0NQnIU2bAfgtK8N4uMDKxFH9gl+c7v4QoIUqmUz2PgFwk87Nj0VK96NFTv+IeFOGgaGVofJAzjfq
khDJNL0tzrPE8NdDobKEWB/jCUCwh+B5gN7n+cqakH1sTcva4CakmdkXU5xKxT31lrtDxFYlbDtY
hdTLM1pgDOTC6FsLAn0V8hDSTv8/W9cSO40DIDt5ji2hfqwo3kN6hB8TElkwk+3kpgK+yHeW/d+4
ABhhAFEAJdsSsqt6RmD5BRP50xwmW4IHPeiipWEuYMotWc4FygQ1ckd537qJELjpKlVtdVBU9GV1
72K83o0iF9P8z/60aJbiciV6/J+fShnjay7eLALjI3TAs9r+HQOGiuzISyNiM1AFL5UiZb2cBcYm
968e8Pv8YSGfniUiKbAOs7vg7OhBW3bCtMduJz8udhYxJG2SfBjXCN81HRTjeEvXf+pAT7AuGMIh
g9NkH6P+t7MeqmOBv+1ahlg60WOBxCjXl4c0r75v6efBiRRCTCsMzCP4pLgkweAh+hthv1yUjgWA
SvJu7TlM7KDUWbiPMB2XKQJkmhkZr1SyD8hL87XKV3asST4GADH5BCY7hoWC80ND5w+zOKjYTE3S
kEHEsD66MrjsupuVK9v59mMckdNWMPmyF9wtpFLf5qWhFjgZP91agJzD69UrSN/H/05Aeo+onGQ3
ZktVJJdNR0r5TDb2ufpsCZxosR7XugZtmJcTBLG80mlh3rnDJ4rjZj/ArL/VzhTiyk8c+1L9rtBo
8XThTL4WeYl6mOi4MItxdy+h8tarCibcQFQCLFoCwksPEz13Rlk1ncDsdL9wxxJZdVIjDpZ9aJJC
OOTq5wEaRrtgqJ1kMJMeTvNy8ZjxSSaRlAiIMENajhJbL7QIttu/DRvsaaFMUCe1v9jnYxIksC5D
JZ5qF0izbZpVscllcJQ6L5h/pv/uJh67S7hWIBrABNX9gU0GUI/My7M/EChMbv9PCwibUMPSOo2Y
vGVQD34rs9+ePgPyIxU14mOqrbnzm8K0APayaJzPXVDml2STCYuvkPVcQU64US7/7QIRLsaJeszG
kqwSIoc4T5o3SZs70pezzSJLtn6w3W90StNZIJeW9Dt4vdueVUEidAEqtNy8RG9668kBmldUoM/i
jdkuEdB9aQlMN11oj23Mj6sXl6KNXjZo5G9cDcouiklk045/JwSZ7VnjOm3HgOo26GtZvILMtqvP
a+kdltxfGNtO4elEH1g6cKeE9/PZClkj9kd+wGXOdIGQXkpeD+ZeuZekDb8MPbSs6T6PRLVCmmnF
BcQy5dicskKwR7GTahM3fXWIolO1tEjMqtkDU31J7Gt6gxAvJNVtFtNHAi4erdzOorhKZJY7fzE0
77hT51OgCetP2/NgMFFo811TN+4hN3fGdNxhaY+htKexevNg/y8AElbMw94DO9VDo5VdBhUs5Y91
LijDRvcHjXiq4FffyxgwhgfPbXwU6JxY5mWbXxVA8x+yiGWh0S2SZjw/eUdi5PjRZCTq0hrcB1iW
CegAZ3FhultSS3rL4xBjw8Nz457/2CUIiU4oe6kKhjDuA7JWDoW0DUvmKZPD9W4YvcfBEmYiaXWJ
AyhLK7y7oX0Mp+aYmMmLqB+R8nol5fEVa+C71zq5lAjIkdxH8Bb1jZVrPcWF4AXoX8cRRmntPGDJ
3W43JcHHjUnok3iIbVzOMShajJvwb2VnSSZVKe960tqMhstHPYDuSQ/gW7jGqBRH4yMDIlG9VCPf
lltWczvoOedwzxpjpHaXfw94OtFpNd5Cj31AnHWNYNoCaxsgCeIbvfniA08x+TUyEBig2r7wvFO1
U4YlISI5/uhB57nHBJUSPrHDiMpetLEf9Lt+Z0uKOQIoQL1WYrMAJvYvHBMsIlJLHgKjMMEX92Nt
OkQqMgAeLWfMlRUXQ4ppZ8pmnsn5ck3wHw+Xqosjeaeei17LC3DybyQHLA+N5VoOt5wz1gHQfVFU
ojAGuC4cHObT0fPaN1KmvviZSBRsFRsxS7RoYhwdT2GHKMDv9y9EYFBxi802MCiT2cqKp2PBHUFD
WXymKKcJzicqzAQIVUxgpoJUd9GJ92ckEVOY9t5mAmc5RBT9Ne8solcAMO60BLYaUzkMB5JAzNwd
sE6dIh/paou3IUISIEGF4K6YxDy/C1dFGl83QyWZUF4Mxzdqaq8RFWP54DBvzZuU3Zfw1RBo1M81
zQmxrYeLGRPBYBckoK+1bxrpHQ8oKaw+Q94OZAWqIOGemenGzdvbxKCqfyAPIr6XKcT6vME7ETI9
c19A5dsExqCwjJuh9J1RdLAqzSvptixfdDt7gwhskBvmyFeh5OLNZKCbvwXuQqQpN5f9HoeYW8h0
lR1bMrCsVhFNViyC9+rIthRZ544mZWis9Pr/zEU5eBex7goO1giA+LCfmUpUnRAPqUtTLvzuUgCl
+qjJ2l1Cc268PNgkwsj+Yt9Mfz/qFMgGbxt9kWDiZ/IfeFS3nG1D9rYJUm9JHnUQZXbZtw8VQj1K
7+zRp/S1BSXkqa6LyPSRUSqH4meH09Ow4CTeyNlocs8PGu++6ORhwEx9t7mKI5t/r1Gkp8B1fmIs
1D2NsiT5sODkCtfMos+xdqHLD3kn2qqeU5m8byAdsB6YRJcDkFpE5lQGrP4GYoJgn7ULyzsdd7dG
RC/cfxPRi9ZqpJ+HVTLv6MPVlfdBiUw7DhQocucEFvwzTZqcfrMER9s5CegglMA2+qadQVEvXhqb
ut/5/A1Im50pNYrpCCeAvkKPQ06XydSf83cfnerBnUgfKEco/f3FnEZMiBq07pNa9ppsNftl/wll
41jNtJO9HeqLygGb1hQ+MMAbfZffEZO9CRyzcXjpRfPwB9Xo3oYVYQt+Puu/c4H6qCH3T4Q/sLqd
7woKBvXx+8hXIt1zTEQFuY4fBPyuwCcxtEB4vvuGAVeERB7KEoP/4hioMKiA143GVtTk9ysTBLAd
J+lnxecLtDmX28jDdNM451BVsZsp0/a7+EWlYv3HPYqm1e4RqQR+HcUb+bRYz24feF/MLg7KkEMY
qRqV5AUgb28Llm2k3qKly2ocVMAXmruRZJjR6BEPTEq9A+VA/dzYhI8fZtiZeSz2yVQu5RhNf/Sg
AVz+aDFmIv08zaIWrTe96U228XfT0ikQ3qCG5rs05Dz4DqCmlymdk2z61r1mvfe/TarWS/ZnUt4s
WsYFU/LxLBvmEjh4i15jjCrg9SbIpa8jHsKTU3H5zCfzGmAgFr5DFiO+szrY5Fttuh9kYGAqOUcH
Yac+PDk1kEfTGib3iwXabFSsz9IVLrI8bbkVxA39qeMO1DDY/9J09ezW4z0ycdxmI1Pqn90ts83i
JHDaKbMOydEQQPwM7iuOd+x1g2/tm0x88BlvD6JG+4bC1OvkagV9nn6+0UOMnbl+of5wuZ6CtgGu
EpoPg4bhsLB02J5+yrWaudfpggsJXDf3NC/Wl7jjTiElJd74JKPAiBumVSH+bY5inlrpbYWpGNha
mJOBXOPVxPI2qdDxKFNQTNCLnvSgb3hHWDL7T1Mwlk4ZcXpcTMNGuaWDdEna4l4NXf/0RPWpR6G0
AkqtJw6ITpfKuEs0EKiJH2jD9IpQ39N/vv+uOEmiWSD0LEBAJ4f5vkdXNGbjh8mde3tO0BPJ8yHK
4qD4CF4GM43a58eMQCrXBKHqDYH/pOhrI72l0dJcTFOehkiFu4VwsujVvCYP4Yj7+Qv63npACmXI
9QinAGy093fnM/iLGx/7noRgIZoV487Ngy8K+4QtwdKdkH1WLR1EF5RZZUYYzrEAgfofalMLO6fH
u6JD3WoiCI4m1U4gqtdlU5pWntQulqY7gjFlLa2wCKt5JvMbxUxpDX/d79DT+9Ogw8K+jm6EQoJJ
jfPUlvvXfYXysEaSzRdwufZyutMctm/i3haep9Tw2OQOh9J7OQxOx2qofydbs4daVm8EVeLdGlg+
T+8YlNprGzcvZViSi2XO34+TtprJ3u1+kUxI3S/kkpbIRViRK2P2GvQNFTHK8SuKCP0ovpXZYO4X
TCYDQtL+oij0h8WogayiN8HknnPqIbav86xomnSc3cFPFkqkk/ZzSoqxbIAgHhCW1QItf4UyYweQ
5FzzFq0UOKTZcZBLl7Vv2byuyPU0rceDqlSzL/fdf71mHsY5/QZ17TbShx3PqXA8byvWZNi8ov9P
jLiGkOuwOFDLwEairyUGfzlHjSAJfF12NLIcoBBxxw/uCgYfgJXb9G6r72zZbt7zK16Z2KA17KMp
XbPIl3F43nRgRYpHyfRYkERtSGtGBgejDY5ZulIgcHAe6J9Tv12UcpsTRbvEfHbpPnztjBGioE/C
PfEPT8I+38cMmeYEgO8UH1NGbHJckWJu9QVMJ/duHxdidFJHHRuWo7Sum8JJSosQrY5Qyx3RXMbw
YIDeFerpebsT6IH4CAJ97hVrU0AfsOy9nfJHGJasB/zS8Mw/1bAlvmldLxHXCwgl8IHgElqUJCZb
JRGLVakyjJWKA9NgGh/wS8QNopIqpw9xBI55a41EaqLI4rljkr6hLqy76lrehyimt/Owb+n9JDDJ
4DkJtZg+CJkEvZeKwW0AwXcx6JBIECBybBToMeUANImEfq7sv9t1mxNO8ZVCkUuhue/wHTPq9Lmk
J43ZB7zeQX7UZaeI/y0PC+/fXQJl3P6+kS9Wngqo5faPe3+db+TPOfB1DR3ZEZgdjhzfdKuV+pR3
SyiZk8e0vYcyyTu453vmtf/UcRbfPcI/CxgqoJBue4J7z8EGSxnqxOEYK9qXdPl3WK1wsmy1RaSW
u3EquWpenFYm+8ksBSHR3WfWRE/PMvdVkCYOJ/zSy2++Y8S6MvY8PsC0XwwI6SytW6GSb+0g9Odv
sEgqEaGBQar9r0JQ2uoMmlZQ27VvrKS2FHHBxTv3DoUIYdeZsQ6ip1ccoTUSVZPSrU2bXCUSTGDO
+vaG4Sdcb3Vx/OW96CqSRIWOzV5zsyxzF5/vemFUQlL9Rykp2KhrgS6nwbkFq+5Amy2dbGv1t2jU
mwzL59E7ulCj5m0f7wABs7EeG1B0z42c7YAdZNyAPI3lyDVf59DIkd8Y6fqqIoqCAlnuvzvPZlNT
TF+9x37b34kMXetW0qpAR26uyM2hXVJrUdHHFuWHWVOnxY28+wuRp+KuOgfp00mvxR60Cb9imlRs
/bb+vvqYpn3/Mwo6xyzlCbuZGWQU6FrMXnzg7iFNqvl8jcVDZm/9WNDHxV7z3S3yvvs9eCjSN1+n
4qFrwpzQm/DbnoNQuXSpN/as1tIpF6PIMB2028Pq+uS0Uw3ao3WJ3Pldznl6CLu3JM/DZLd/snwu
aVpk/MYaUdOe7GdLW63lxFRbe62OfUUlmI4bqa5dfVKLt80W3Trj0yqEeJEyPdJXyy6mfM6i92Je
04oP4QlqhAp7w1A/iNZG6w8B8l6pAnVir3mniJbzGXF3N5RxcSI4ZoFNkcpCPhzJyJNfnhI5uNs3
PMYtBOPO5hUKfF53lOb28pH7lRvgM5jYP+WhS/dA/quKBj2wwF6w3gde2Gxh50JxVv4r3dEZgyEk
ZFqkMB4X0QNAkus7x47Y24U2VGOiicalW6MR+z+6aAmvPViEQM0Swto4gn7viy5iwkfQMSR+piVz
0qHLObY+u7va2aYZSevblCkerhVjc4fiaCYaRas4oba3r9vRM/lsb/Fsw6OslokL1iJti0WLHx+E
BJIE1DCRY3Iu6K8ECzeGRdrougwBdIb00cRSi1lzVnunpiAZkyltb+oHrro/hhrk/d8jWw2jSjgm
1E1PLkw1MNBxMfNslqcRxEB41Y5vE21Oe65PWTdJnaEngxL/fMT7YlQBHUSnzxGLpyCii+FPX+BV
UFs3U+5sUyYHYsn5Za6CmfJdvMyuwrIZvkcmgVyfXe7D9VukNY258XCvKm1s5Oib6jTSUlyxJf+D
ZPwWxubJaWEsQe26xki3X9bm+pXBZ9vQEXEZQEmilhwTIXB8NDSrWE84uwOuVmJPnB7Kgce/eAEm
9XdjEr2CQ7JZzlNv1zlAMANm6a7vnTshK8SH1BOaNLA0NYaE2TNGDWGe8I5BgZF0NoF6s7Bt57AM
JMIP6e63IqwGvxDk9DCOkDdK5k4HjRqrJwQ1rJcZBI5SQSWhD/XlfBq5xfIXBu9clKfJ3qiDm4V3
I8wSPigVwRO8sCsIQMl4Ibktx/Imh808oP4wUC9V532dQTYdi12S9RHB9iE5uokoXAQM3tweLn2X
7S7ggozJdk0MnTdpBnM+ieFD9s5HzGY7VKGBe8bz76FBEzlfPxi7GwhF0sWUQdu+RkLwEGvNG/sB
159xiIq0hciENnMyMBvNjXsGvbp/SkExoKdnvTng+WzSMavwWVAAhr+qtgN9dvHfljtdHSEFCjLx
p8upxwHiTvqyYbbXdJKpyHvCGXjl3DG2xTu5uaVchWVemgutiCiZ0XLRR+LlqZasgnI6fq/L4ppr
3okpRJk7TfMKVHfAcHsg0yNm/F4KtCCLH0D9a2xvF3Xtv8zGQqaltIy77ATlv2Vp3YxlkuAGcJmc
lKeW6XybIjZZ1f++qP9uVAO+w8nEUyH8MgtemhKtMZp4Mvj2BstTA9JRGqzCsH05qP9WDbsZWxkD
Ilc2vA+XQBOCWowGoPzqr+zPGWHJvwrEBXX9IWHnkJ84jwWVoLX3gIjP3HpNubG9MpUHW4bTWTod
mP5r3WVt0MZ+UR8qS2BlqUYPNp/3mEfxMrFKYgVjoBneUUAfcoo5Bncpuk4xToqEiVecxC5+k87I
7zyP8o/JJZNzmol1P4JVwtPVGFT4MmtgMQp3dBvBH8kp858oI/5ICjKELRKB0YGuCWtZ+ZpIUupr
WZ6TrtxilW3B7jqYxrYisltcPPk/Epav3l3iML5NA9vzKR2Aa90p+HVb0NcBTauMudKRh+oj32SX
w6SdA430unZEdLAr6bTVFsL9vDRhX4ssPjkOcR9ii2iWHJBIBO1oeqAfZWL5uf8DKk9VBuUjZKBL
ffllCr5YmeKHiQZpzg+fE2SoqT65pqcDAyYDkJjDcsHnaGAxfq4XVqSAfSTp9pcZa802UoAcxbv5
liHgH5OFhtSFUupEgH7JAh5rAXSTkb/MD4YQT7gmWqHoyMjqZ2od0AB/yVluMT8dHnh+NpVyiXTS
b+F+THljToZZhK34f7ZtF7VzMneHht/bVNebBdjUbH4Q1X/xqpGzDpGweeEJ3P3EHdth07RnzZ5R
Jjn/KLT6UEabauAelDcSvhlmKyO5Vbk26d0ZJoDSZ0UESwB8wC0LM/02n0jWvqu359kISj9zCuIB
aUuT2Yly481Vu04/esdM57Y3He2CBYommb5XEVjf+MR1acrOCsM2r4lnNQs1EfT8MAx8N6gANZtm
9TmAiJ+RXgHa3faR/BiDIO9Pulc6XTctaetVdD4g9b5N8sRvlx3YebdS0NmUFgTjCZ61sAq7zXax
jBXrc3pHHsu9zLROXVHPYcaJ0WIQErZpswRq9misCgTNNm8phrbISatewdZCZeu5TkR1o11riMLD
37Se1QqP2/Uku02f7HW7p+W5BN7tIuVkJOkGPjMXCQMxWAG9butXXtosnJ3g4XZ3Vik9GE0lTEoJ
YFm/MEdaUkpOKNbU09HuYu0gFJw7wQxDiTpbtqenbpSoFkSzd/lK7styBJwp2wEaLBtwp8e8hJy7
wEHPojICA5MEkOkJG9cOb5+HkmrS8kCUXNFZ1kQ1FAdlUNv4ZAfmzUT5AXGjqzU1tmTX35XlPgdE
xeWHTWkheGIcZQAGk8ArQVNCLMZ2SxYv7csPgJWJriokxnE7WI/bKqd7jT/DpiWL37AV2+fmRZGe
221mmO2ZIlX0Zz5DU+r9g6QK9GYipC0wv77wfv2cktfu9pfbwif+LwedKEgKKymxnjkQ2lCw3pkH
HGU+vIh/xBqZ/XzlfPXbOupSWjNL/sJyarR3nP3ZP07zur0vQH2DXUxbE+k7LhkZobOYujcjYJxr
VC5BnuXVzTh50NeRL3TA98OtAPhI5Y4NhQJf+5dPDAEd/hmIKqMWIjGFNm9IiK70HK8AXckbwWI7
MC9ZH32OgHSZmGrFPRWyHi/cPgz6ib2Vwn36eZp3lcu/uu9PfXTQafhimArOvLHj2XKCLrIL6DlE
wyagpvMZgO8/9urXQaVJzZOS4hxa8jDIMBd+7oO/7K7v4LxEAKoqoUsoRXDQ87AWhpGvi8CTfwPI
WgjSIAU4IBh0wJd7J+EdlqU9MAg7Cy1/d6xV6OiH63zUXB093U6CTWza0S+ZYJHZPu6o+eu1QG27
v4PWC33Ia2hBzdPaUFKxwckrsqp5JftnetiMjKOEdW4caet8sAmok3FqkwKfOoLH4Q3IjgP25hx4
WHhLYTR2rl3/fHFgLpABGpEwCRgaJ6bcxWuN/B/6RXGoRQhATvL+hDSD2phTzl/tiQ4FDbWg9R32
GfRkL6Xh4wNXEnG+ocSOD4A1XI5Rq7szeXDiIEc2cZb/f2oS+vmgFNcmbMDegwsujfFCOzvG44e9
AXMnoYGftg4/DUMj5MgcNh3kxfKeG9Ukb6+bdha94AXeLD/Ct9DHUOLwEPgmXxH/B652uUr86Fwm
PI9UCcrqRIV988Wxu7hZ/TXtLJ4tUNEgYcDSl2bhwhsNoHFovrLe69cHCB28GzSbKC6xu4qOf+b7
bkyDR9vBuhKBcR9m81j2LaPfQDZIJv65wVmK5hVTiOwWwA1+x5x2nEpu+gEwvYQN/pRGehJox67k
0YIlmAbrRZakz3v1Oxv3frf2zn2haaPmXaulmTzfVCszVOxrnkklJilUXEByTLSubE+uAWFviWAL
zFQALERLP3x6p0kEwQPADsVGBYVreZZNG81gKuHJQWUWnSwYve0uV8N2uE+nuzsMOxiXuWuSInkC
wt0vwJvdWnXbdkUkzmn1ph4mC3RJcnF+vV/2QSiYWl50PuA1ML4r9lRxl5e1E2LZTDMFdoWWH4DP
Vx65jw+y5TJ2/3Jgpt1CwL+qlrSdrd3gXQKbZk8jMN9YxYOgak0JvBXfjGwvD8F6sLz4ixZG8gS0
NiK+GOICFwGmgmhqb33fzop8PvKmvPttnKWDNtTy3x89R3faLVEZhpDcao3hMKO9+pKObKffHYHX
X5+eEkmask2rB88uRCn5QtJGNLpkWuilxiw3I/k8JI6rWZaf8SNsa4zu9VQ0EEtJmk4/JmQJ3kO4
Os1fFs8fk72GYxPZgtDVb5f9LatYQpIcQukbyG8algPbVoTLMJkukpLh1d1gwV036+JGxQMcGA1O
7rFDyx7c8zpbdWyUOID+uM5mtD1Z6bnjag30XojKz/5+65t9s4Qsoq4fN6Pgze9qRQKCusVRf5KS
9VEFP2PF1Tkjockh5Ds0NtRXJhyeBX6Tiyuu0PCVNIWk+zzolJtALYUpNvXGLlNMx+r6xyLVQNTr
RceZTaOEZdxdN/3ecBFV0n9PGs9MTazVLffECi36i+nlHHWmRKs8RuYmmkDYCL+D2y4IkNQRbpKK
vCq8tR4J/PVW/0lk6ZsTMiGZLeYOBGGdLwmiiAGjf1GYuZiXnE2D0x5d58APEpkpJ06SqVZPGwzp
4An5qX129iQ7zyZIZFXFHmzBMZOc7sRSNmXfLLQqg/arBfMWd5DX16BdPjdAkPF8psrAvfC03m1r
eqog35lgSD3Qky4ZtlDq4lRzaqQ6MEQZhiutZ7RxbXUZDkAHEo3QFOzSUxIDlqwnC/u0jSvoaQBV
O52oEP3oMAkeVbHZBVgK6vd2Wh4a1WVeKY7/ErK6L6pSaJE1u/rFXjBNotCPm4lPOkrRZ9B0D0gF
V10miH+J4cgSRCY9HOK2D3bEUGLXF4MmUbo323m3SDZv6f9QttGCacw+yp07X0mh73wX2Tn6+u3T
sQtG0qHpsHkwddH9ej6eTMGZEjS2NlasNsMjKDsRVSlEMU9cnm0h1j3S2eqUMD2WhtjdnYWANocs
1i+/iMA1X0eqDb7i4ihJ5K3BHM8beS9Xohql2w3bRLlpQGan4ObEdYE9EPMBi9qHgZAhZo9DW7QO
ZVY3XCaEf/udPAyofaEoT1FMreHpANdQE8BIaUx9UvA6wGrceBe1x0Pk3G+MyL/HAHAH683TACpL
7aj9HLQn5XLqCaFlTAOq0Y885ah5vnuSByfjMq3BKiokldrqT9HZEeIeTWdk71by4YBElop/s7Um
vhkULB9RVIRJmwhJzt4Cf5UM/Awnoq7S1q50C/QMJUZyq11Nmq89QJCu2vWoZRsSHBb5+9s2XoXV
OhhlWd3gHd8/j51Cu/HS8TkKBJQk6kXYBiZv3IQg+Dyr6kQlNhdBxcJsm/zTkPgApNoLuSwWawcQ
cH+IA/r1VhW8+st+oEeup8in4wfl4IHH9QhV1to2Zti0cCGJSqQNbqHRCFd0Znatx+SLgrkFPZi/
LK5Q6Z9qvUCwuikGYUse3N9bZ/ed41uk/Ne5+YYDHob59BJmPF/1bRON0ZvtTnGhbKnx1NA6WXkG
T0II7pHjYEre9GP8q/871kLhbne7lYzzHygQxj55jnbZnVbeqelEYAaOpYv1xB49JcoFweTZuddt
PGThDAEtZKNlCLDzNvzHet66ObqPOItuSwa5J1NMjFHqRJLcVIAS55l1eUjua7BqgosUh1BncKbz
R3kdGHVN3VIcl/GJW/hM2ooMuDo+u0dUISoeJibIP216EZkE2ImecLpWINsLnGGqkdi5wFSbiBM1
GEa8VP/UnHQnfSHdIYoIt0LdvvMvZIXpuyErKiXghO0YlPfZlHTwX/nGKaZW+Y9caOfsO19PL9j1
IunAaTZiiTgkXDXZOMSHfeqXXaSCNQ78F80hXtmTW/PHMBXvjqJLXAbhDoUNF4aVA9lQTKNC2xI5
hHediLf5D7/kGN9QSdm6B1GqSSkHR8LR2e1uZsqksoil4koUmXJ8fFmB4Yfs9n6bZcDTMsgqhR9F
zDbJheBEKCOmaVzEgE/EQZZQR+/9H8v3hgb0YL9w+qB2xfv1VFfmAhDGYTKYr7CyWMC4HLEQUh+7
ALbNcjcVZn/TA4pDbh2Fw2pS9k3XqowtmFhFHjHHSFTKJ5H3k0x1dxuJzBQkERUb+g0CpeaNvszw
yFwdF66g4qbd+3Nulqip6FE/q9s+AprJmpuFzCRszo0aBlM6hR0OuIU/2qzb1be4PMjaLeQVSnYl
TvaFv4B/ygCLugryhk+Ef/Pl2mPAjnt7ATq3CE+4O4wgB9D+bi6sP82HzakbswxGDApy9YW1gVg8
AvH+LFwUa9Cb6ev9XkDgBenlxRHb2T628xeF0kremIOaiS4E9QqOlPsvI6QaSqLZrMEC8mZ6MzEm
kQY5q5Au+oCUiWPopGSfEilWJoLrKjlsR3piLRO9Rq3z4EuD/ZdsrCLXxXVXr3gt/vauuCoP0wHA
c0Wgvdstekv8rTf524JkCgSLhZNUj5mY796rZIgJEsuavgOlOtWZwLokLQtVzCKAUyQnEsFLIX0H
7hOkf+v+kyreq8HLggHCB2SrME46JvGveuSHaoZhHtWb4smTyt83cE19A8rgJsPVhHVNhPuL5W+5
zzE/dYLe0ayjiJhrCNmWxEh2ZXm32e5mIStxufKnB5sq31J5jJopo+gnSsPtqe3xpqKQqiYkYdQE
QydS6c5jUQNhMltllCftY1iIFFfTM8Z6X1Lbat07xdVY8zPgrVqqjHaCRsNtMfRFafDvbW7/YUMH
Hwrh+XC1Tx9X+hwKFNIztJJFzXgGKQC4yfKcFy0F1aaHaFuKHA391oAl6iUq8hbE5rrnhZwsLeBH
aHsjjn+21HG7rxxtnw4vNS8RBJ6WsVJzPOso0HWRVRvyG92C1dyrqCAUbERyUoN10ygcVqVQ4ysI
8PwZrmahfzd7fRc/J6oHEkGSBJdVXtVQctfvME66MZ17s91xVGtD3ozKgnwGl+bQ0fX510pbSGGS
slUcOvCd01FrmoH6+u+4JRJ+CJPDJ5BCDuSzGmvwjsm1CdWmx+QYkx4q3fpbogcD2rdztLisTU3n
W0PeBDvTAKRZjVonRTeL0wZK4yAzIrBOORVblYCPI8OQQWlcYj9V1td3DGxMqhoAp5dsOLcJinhF
3Gz40TXJ+p1UwJTe3YXLnFNNeMmlCrpXe1itd/9IOJVylPOeTqccciqLv0bH3DD5E925WMb3h6hu
oeL2wFOcqoKjPwmYkRXM93G616MpC9KsBMvSQ/ptdh9Vcx6CQySlOOq1ozOEX7RcptiTid1TuX4d
SLxTsE13EdD5QYY3ML9vCe+E9PhSPuwXXq/6cFqcV/AwEXd70jfk/96oIsyaOpvIPkNI+KCVeXFX
DJv3NGbWHc4tw7Wgm9zZBeO1zU3m4+LF+Z79RWLgv8w6aFdixMEpOB5y08stmEnbb70voouEuT9X
vbJU6jAXHS8UJi/Gvm3dzHfPiCp32NLwION9DzCzgo/GdJ0EJkQs/G0KiPdO+gRFltjuVnZaw9FR
VridKJ3jV/2VBZDI1V7L5l829XoDidA3NMp2n9KO9ZveLsW6MQ+ZRtNUcNohWVYO5DyaP+SxkVPC
Fn/gcMlk5yn3sx3FQZP2/n5z+hd0NByTq2T4Y3uS0MoaBrMjZfafrAekDA86uL9GD/VZsmTcVQY1
uuZtpqK2g2i4O9efeCqdc2fe1SgH8f9O/mwbsjpFKwohLfv7ufdo8BCnnJOxbij8JXX/jyIHKQLw
l3W0mjzi6utr6y8ImlXjPtL4/kh5fHoZCex+ZuAFQoZktCDM5FvJUrt7Hhy9WSOFHIeJ6lL2lXFv
85ciPNT1BBGcyOxAWFcejf1lO2YfVrLYLuvoJ4aw/mrdqzNvFywYKxOR0TMb4qQS6gGLWGlMwSJI
3WpfgK/vw8u5G/WXo3WkrqFO1Nvu+IQ28TEAHXARZsSbIWgNR6zOK4wXBZK3my1wF+tibYatRr83
0LE3dq5dpU32hYHNSUaYeIr1UWmmfnccmQaQge1uagP3MrPx8nKGXk7aFDYY3HQxlUnaDHd7qOVx
btvzP1t28lIBEHwsryt9sy8ZNVklhwEkXh5IgmmPgfT3w5o232G4uvghv0CKpNBcdbJpLCSI96TB
pfMTxtN1Oy8a6pMs30LVjb8OBxOIsicyUYCb+s58Ql6hnNFwV+Dg2DlS0K5SKYdcuCORrBngPwrN
h5G3JTBPEGtfReiruAOyIgDArFasAucTn+/BWlk4b12o4uVVim42JjDhKUgqPx7pXFT8wAaeNSz7
TgkTljBCF/pGfePOCACgFtX/WdOp02oMCKhQVAQCpAkIIkzc9xS3NQUqEz1RvCyjt+XH740Ymyfb
75yZtaDzLZiCh1rBF1KK4m7d7QNYDwJkPfdX/NF95QsY4kv4VjTpcgNi7Fg+x5xa+Z3/jhgJjCK6
/9L5Iuhzo3oPcRoliLc3s6M6KxlR/9os5RvrOiU8M8HxoYabCbxSM4oBQcsFM5/JU9D15kk9KUYs
YUDIl44oRsl7aCioJERK8TrN6uk3PJU5RX329qq4up/59b9oMM8AB6667YXC+ChGJ0xLhx+vUJzL
P4Z2LxNtvo+22iRGhiy8HHFW8o0Ul+ZlnYXslHQ3ZxL4G9QWCKDyI1D+ichfQ2Bpx2eKpOpR0Bt8
hwGlz+Cp7r9b0np+oHVI8yr3VbP0ZtHWoOicgMM8+YfmBnzTdziMz6i7GxpY+EB+gvQhrCSttnUp
/Q62Cs59t5rSt0H21DKRB3RlMGbzTfH4WgSsnKdF0vSY4Z4FR/jv4OEBsvcj4ZWZF3fvIUxkoh2D
LCtDcSGN/rOzHLnAmB2gkagFxEDAF0NcFhUhU5wLPvI7wbGgA/tCplvYU/EZlt6Sf/eiH6vYsWcE
rHfUSb5ooA3SLqtXXmG9WTBize5UCIFfsi42qRFkj7+hB28T+bJmrpM8ktgxIZ27ht/TA3WJA2zW
F50ywHdNf+o+9honaLdW6ffcVYPkyR8vcbTS0ib2Hi0R0TCSlZHFs77sHk61Fyo0kNpr8z6bCTyo
CIDolJXSsaGrNDZbNVxqo5NOl0bEYFWPOpptNw+S5ht6WJtdLAEuYb1QaR+RRyW8jufzRy5ZlPN7
ItpLk7pLWBouCNN6ZWGaMC8DPLx8rgqsMfmc5rnTTLqHGKhqntu2u5vpnhlMakkTOGCEDlqLDTdq
N4Vf51m40cv7NDwpE64ZavFvPV6dQEaOSsReXyBYM+uwrQPhNvllQNtkDi89dmYLKxrZNyixz62o
1b5smvInWq7NCCDxaMYrJ2DNkNY/OexB5mDkqWKPP8I8ecoyGcb+1oojUGXx/PwiOQuSoHriPYVy
exQbyW1NKonrt2beoptOdJe8Kzfo0f8f6LFMdWVM6AoeybFTmIDVm9uZfXuyxeAZuFnJATP0FlCP
0/te2DKHr7lJ0l2Ox+OiFCAAtGx+B47ibSXNHWWLB5S2gg6tPiC+T/0TMV7QzTLVUBi6tBBdOHnK
zorxw6UUKvcfVcKQ2JzAf1x0wyXRrUwU1sS+c33gorfj4baqyptJmNRZ5/dLAj4VlmQqijsDFBKe
D9US5nw0GPGkNH2uG2GKJbzCcKASFoNNOq3iCYZuuLpFGg+KMxjgZ7ataZoWpFqEHLn07W/C05Yc
p7iYrZTT/w5JoaSmjOhlF/gWQa/YWMZ7Kwcq9xdhUwRuaFhAO/FfHLIZY/McLYUxVLIkNpQN9t6M
e2q80BfgofJZEIcQML/zAb889sNJTP0hfjMrYIWCUvz4mAOaaiXHxfFXxhrHxxplQkzfszkJKXXE
V7d6wsYobX4k4ahdnfIuoUyYyuc/0GZ8feUustoxwpZMZx5udcYBWvoyW7kgIc2THccxsg5GGF+U
FolTH07s+dVgyB82plQ4JEGJwsWNKAMSPWqYpTohz3x9Qj0SsXcSv9gxNdpbkUlhBk3H/MeAqHtS
QObOwseAwhwDZ9pppeaKm4452yHIqizcR7gFiKU4Lddz+wuODbIncmtJmN8vmbNzWrJimYQaSMBx
qZoAPrm7tA+vK4JXwAGWuSF9MOimjWgiLW+HK/Cxl4DwmX20JySjXZKTjHpn1FQmdXgSP4gzMdO+
5lYwoLnG7PvrPEmbVhTb1ZoRY1qKZ3XIoI5I4ypRh/MOj6PW7ZHKNEdHl2dsrRFofbG+D0hiUrd+
OXrwQRZ6ZWSm0hnsTv/LlaPuq8Gos6yTZEXTfAQhHeB+THXQ89G5mWRHqMqrYavAT3c2k0o2Zl0+
L0Bu3CbsOvdg7ydWKIm1C5ceNybLAExFskuuVhUwDHtTO8CHJ8s9MeWGdRpr32SlSaUSGpPRevx6
Qjbt2BOrMLpiPDuRzK4oC4CwKBXsGZjJep+oO7hIaO3qL8F436mYQTQxQHgVfEEOxZV4iwrDndR9
OL+PZG6/LQGg6mVeffo8uFFlyBJ+VJ6ML3l9OjjHHFtERzF2y36vIoExhB4ppoc0lvzCkRyBi1q8
e7NkkNMENmbZgnAXzuUA3eGTZrQ8zWqe4DCPvWoXPJy4lZY5F73sP5PnmUwnzqsFNcs2rl9wSYps
aRy7G8bDzqmeGJlimn13gMIOMlId01b6hnrNswrNuvG4vE2w9wHvrSb/BBpLD4w+S5np/Jd5dcsf
a2pP8nqczcpWeu4Ivy4qWeBsamlOuuy9pa9Yq5FbqMIO6DWnkqCXN7O8VYkS7ysrG9LMRw6AD+d4
jGWhzpMq2iW1ydxKMAVIXG99t0Xct600dBiM7KXN+Vn0mT8uMI1+2I4lAP4gGjZZ1KicbhMydQhN
rEaiZUuSjPFej12Wj9Lh51/fMZFU8EznhmBxMl3a3Xe77TI5M9bR+dY4NWPsQs1npa+3rRFzBqu/
vDoYi+w53GlOvH3VNr58mr3JsPTGlZL/kCgdUFxIf9S4Pj1Q6a4i3c66MU+DS0rGXwGjteKvFhGT
eum04Dt9XWUJXZ4OrHGF9+sUVYoTQT2Xo2iCMgp/Xh52sxBPahIloxyfGXWGxeReNiwYwMsBOn0R
YUr6Co8SBcHlThBtUIoMSO012oM1HkXMR98l8NPe+9g5EyWWVWjiezP4W836nsxRw805qX8+4Ik+
QN2BDkuYTkA4mTxF12OoXpX0KFnLfimvjkfeKrP17y7vH8wSEGuUMtB9UtTARusfmuMNcDUbRhzE
OMId/Gl7NoyEq7ESFirYxbdaMkxRTyKhjWukbPnDbhItU4fxc6VThemPgTGr4NsDA9f3wuzua5Sk
XmiWglE5M/W0Y4WEoVAo/biaAYnCMOEPgHznZ1bsMfVXI+guejR/JkjQJD6KC0bTZrg9xI0aZds9
0JNdRUQXU8ANEZcwOmboK3rXHRtebu5FvnRAdpWrEyU90BFPsUzk2iQxxQYHMqKALCbiIrBYyKPc
XEwPCJYQxCexIA/e/TBi9rBDbqdUJwI+dwzugMOH9LGVIIt44buEUynQ+CVpj8RJbOlt+etkba40
cPuAnjR2iRQhRCDbHo45eOwiaq/lN6GCD5tjxwmG07yRen/W/1Ns8k7e2GOS52F4YbxNudheuNlL
C8+ndj5FbJLVPl9ehIpkOf6bV7bHDIEvCKNOQdUa1pONqLPupP9AdR4MkWXESEGQmkVCuMt4yUNn
JUFclXU+Hlv8ba25Ispb6UeLD77mu4kIxAuKGxQBFQjF22ZowBAtdXiVhXp5QX1iKc5ZtjiWe5eW
JYXx6QGJcs6mtkkcRiaPOITx7e66s0i0KXZ1SiKoRCq5sxibifhL2MvIgvlUtRvuX1aligl90eEF
AkO5+Uk0rfnA9p4783Wcwlq3uuDhpSOHs9N2uyAbs15CGgbTuKadbCT7NeEFK+fw6bwghCOmZl2L
ec/Zt3mlOgoGpsU+69YV4VxVtxvY9GVb6ja5ThVZQgWYGyVNObLWmxyH4TJHCHrZjcx/OodoJh4P
OFZ/iFmixVrxjJfbogBn9eYu/Mc77QA76/ZzwGBXoJA1GsZ4xeRxFAilAqaApgYyt/O39rNOFMzg
5qdTzESgeAfstQroXQcb5IM/XESaWKv0mbPTVyutrGRB9iqRpEZj8zjsfHXTtNCDQU1GAtAv15Os
r4add1txCQerzwuCooDzKizFGdjIQzRs1ePfqHwxHXahrH2g3QAr5hf75JPM8t7ElY1jjHu0Zr3S
w+FMXTiT0zo01PR5G2Wb8k4hnI2c70/33qn/bGh2bFEJ3tSVNVVCkevxihaYMaBt+sci4QrzCKyx
ONFr/t1oLRUCR5/jWBNCGNna2QIo5ZDs+a7xqaOOxVTc5SjXshk8xIr6sRJH9YLhsM34rb565VdN
at9mY8XkJhRmpErsXzFxk2+7hFbjCo9He4tRo74GYzadMNA7xMhe8FidRWz/5boTqX13+hiHPG8V
srbgJrSX7nWmQR/75UGNfsQhPE+tfr9B/vzQrWZci+vnckc2PNv6aNBCqyscUhWufuEZ5wwvxlwB
VBFofK6I/MpEl42G6AVZaGxVMEocO26NyT4C2NX0v3nHFvUBc5kuqThBtmv31LPFPp6eIRzBuow7
Y269oru4lgcSElGgegN5u8ze1ih4wp2gUBgRw8riAFtwsX6Gqf6KEc4XkZjIED635z6MbT6e0Irv
buzkAIvC+Tlrh/nu6bkPAKVUiMNGE6dPm3zzzTD4s+Is2qCR4DuRaJ7hmnEgcj5ynf6X2hhcff0k
iB7KxrpqBC/R1iXoL9lu/WzidovJyB1pZKAjDczZupKbYQKIn35/YHpveKGPEi7RVQhnHAL8ImYN
NRQd5SRXd0fhSIUTaNZr2+kczE2w3MUxde6OwEfgpV2AAqWzc7HG5WyOTnDUkXRh7w67sqJdfytn
q3i62scsT7CxNe9A7+bUTdcAmByZIBdOBAXtm8tdEeEXAYpFAxI60zFjH9dE5iyRYJkTcWoaBSaz
L17KOhlxWS1pSabv6HhQ6Q9UpYbXHho/+SQely+6LgG5SrabjujkQSqxEKoX4OMqSbwjLgv+3aog
h+n7Wm0vpvXoLBb6d41KtI9CBb3d6OaAQSc8KTnJN/IkFEnRMWxtpyEllH6h8dlLLMtVtKwKw+LW
w80V7KrVLBxhVL1DfgzDzcEPWzAPFLBOCXZzXuhNJFrlx9O/DmbNqFNR7PYi4TyEdSOONwjbuQLD
UG3uINcIzfc9pBRPmkg9nWMRLOejo0U0Mm5jyirFpkjKo9mTDfHl5naawBP9NJyEPB56mF664Sij
Wnn3Hrn2T+afDeS3TLo9DOh/U5fMdCCzktabrfFCe/DwH5fUMJkWrvlb1ePwTvzBG2N90TKtOkzH
Z4cHt4oSidavl/E4N7MVX2/34YjTGHw8TiM/6+gpaoSujWDv8gCxItLXsZaeMrMYw8menUnUycCz
edIz8iBo4PfuSH5SvNFEzzRkYKQ+c088oFiHB/q68/1gtnF10R+LT+WoKSGfygPynUdhbYt3EoZA
N6hPYd60PSGe30FNbmlBYWs0SEMuLCDUFe4w8MKWrdkaftQ6MKWkTisH5ivQtPQP99weq3W5tOkW
lG3xmIywAjKEJfaEEHURC7t/sdzDY9UCjKqxiUyev5lFop0wUOa7ddKZziIMmfZzxgd1gl11Szdq
WSYW286VkQ8/p1mibOglgYSVa+NLvlB7I1C9jSbFxLQ/ts0cEa+qvbv2m4QWhvrAd4H+PM/iMywZ
XphCoaEN3YF53Q2robocn6IJcSBq4fccewdBYTjBwEmO6ioFkwdZqFt/soDohqMrtwDx3pn/0SXF
2puXbrPZkoNhsKPcxGV5EnM6e+VL3FZNjC+pRSTJos4iDACD86E3XyGekb/kQMoZKk5DYctEmFlE
ekSZHN7lMJ0v3HqnTc8g2mm886CTUbnjVaeISFi3Z8Syku+7gltlzrp2ZWbB7l145Cnb2BGhtdDT
YWbhtiU8Ba6ZN2rITKfJle5jIVbzni2wvSOZRCdVcb6ShGTMdVIPedzW9A0bNKXsWnN0geFhtFiU
/sPu3QahprEs5bmcYTdkuOLQUfGuzL3+4mchBEqqbU9ZAudRHS9LY+a8MZ9eKXZ780kTMLEyCyu9
U5ai8jJC9Jkxl/461SnJ4TVXAVtipV7ycm+Qfooz1teNMCZeuffQpgeRU54Yz7OyZrs8ZCM9fMyf
19EsBaYLdaxG0RnZfrGzrSL38sQvuf6n/0uytSVy8BcSEPWv/u9XvFQb3bOXxxUVMhV4S3FZEdww
D8X3MK1j27wpdbAveS52xSQSNitGrrURF33eof/uI/eTKk1SIkP+fav8TCK/Ccp+oOuSn5+S44dz
7qM95psRyQrwtzSrBjoYCiT1qxuKzyYcZkTCqtLrmZee+gB0GQ7sBO+Sxl+mDy05zybJLEdoST+S
HUwhW2Dy8K4igZBdS3HvCE7+fINwHL/EBs+hurYpaRypoAxdUbYypVpaq1F9eNfGXnmNp6qWYCiL
KD3jPoy6bTw/ItvXJNRvk+F56SsQHPgdF1tNKjnLGoYl6uKUnRtT/K2EWnQKTqkNcu6FYLMmuMGm
drMC8CwUvcy2LOtK0/5oJ88N8Db63aXWTkE51BKxvAOolFUa/+8RC4RW/GbrAu6F2lyBOqXrzx1J
W3ITF3v8cS1M75t32TncgzfYO0w6r57Qlpp98UamU9TCMSzhFMxRfulSP7bUxzpG0Ec4IJx+kb4f
f7Mei9PaOpOrcpgMQ5GKrsPIAh4IzmfI9sEvZZH0riZXRPtkG7P33ATtLD75gUonkkKBYxOfi8P5
uIcg+LqN+dbGRVpM0Z8ZZjy4Y3vXLxjA/Qph4+ItDpeMqY5cCvfLJIXG1e5Ler3KzjW9dOYl1UUa
Va6GRCFKJDB8nnybPc6+7RjzRkIB3kFbac13zalNYGqVr5Wzj46C+gT0Ze90ihoIjyzEp90Ea6qc
KMaF07UUwVW43nP1JyxhkAnuf+2N5VT9qPdABNT6mf2CAMFQKqLL+RhGIYft1N96M0CZ4X5hd2ME
yEiboX8YC9fj2WN4ppGZffOl+dT1Q5YMWRg/0SjDJw6lMYAHYKfJ8O+SKRayrFtw8uCbqZLsUNqd
VEk3qmDYO9LGOrqtvB4cvUPFcLwpEqV4TGJP5CAdCwoV9X0Tcb2w1ixlo8IF8rJeI0WpAkAoHQ2N
dlgDrZ7ycdCC/YTOjtY0bk7i05jUKPbJYfE1TXI66ufVaW2UWCxDk9SyzvHtTAiHmF22jMgJhF/b
7TYHaz7qb5HkvrPO1tco4UW4vRGinmuBeMTgsoEhcfD4s8x8y2aCE3AollLAdYxYL9wmm65s60Yt
xTpUKIlYEl+Dref1NjgGIypb58KGUxQfcVjiRR/WxyNaBxXvxs66zc9ecn+qSLIWeLpeqPnh4RAE
iPWIYq6gxDqGbP9KBT/ey4jJZecS8yovudr9NPA9tGqbq091JlEUarILQrTCsgb2pfefPINw/PcT
S1mj7CNBoItQAv1Bv/lDUw4Z8H6YZQOoQhKfJ/a9mw5jYxSB3vOZthg1Z1Ea+Ng+tRKMawLZ9hio
gBI7hqd4SKFEvMqBVSKJ7f2ywhJWo6lv6wnrrlhdy3RlQTWULkK2Ulu59dAVNQCJadRwLYU1cQgw
/F6LuQ1NMgL1aegAl0trGr87ufV41hY/AHLMxA5kZxZN4QP8LRFz26Txn77MLmp4I58X7asEEhbf
yFGuZ2nA+/Kcmvw1Ytb54JjsNHCl3wLPZbxgLby2/34ZfK2nte5idsFiisuRsb5YdpYSzizzQUGk
zWesv7bJfYu7HB5c9xZiuRg+LASBSGZXb3yYFR1HnrXqtXtBdA0U3TakLP9vIfkRXiriGvnRmHp6
1VU+DFV+aH9ZSKUUSjNo6UXSKNcY1JXTHWdS97vradRw5cJzx0RD0oD1GqklTbkX6nR/WZsTLyAl
aToMAS2aopkuy7NsS9sWZ5SfZCyLbsqgsL/f554HFkYSREtDYzgksa7Y8aNO1K2NsuKY2wfmlpYw
LzHbY/tiUbtcqnbVJZQcdryrJxoEJ/Bkab1kS5WSENauO/TFszF0OZ0Fg78em5+gJUtMAwOv0qox
3VpwHXrqs+AsISf+6T18VZA+0kkNgLyroNytAb8NDrlbbDPMKkBNVQsXLlrN55Q27r2lv3vb7z1n
iIpoob6qKyMr6lMiJ5QQBkqmce83wc89c76f0zvNxsoUZckJcUV5OEQZEbajZ7U7O6mWbDR5ShKi
wVtGVk+S25lf0qfshuzxNFCrJG1ZoYUzmexkGjwixEI8TaSe/irBIbRdjn6LLTdWt15OToJrvjIM
4kCTrhd/HgXNW868JoSnsxjy4BxLl51Obg/eSNGwHwwrLBpLZxQMH0PH+WYJGSQTAtm1N/Xn9eEX
IztAoRayVCkutDeOeYDAq6nGhVIxk/HIiqLxOBZrf/52rbMLu1/sjQ2dDtGLrLpKrn0YrXKvSvKf
4cIxVIhB+Gk3w8cazXKKgs/ZFrWyChpBYW+vRx5P6BRtZEWBM2JBMzVpoWtPWUkC2ALmsHvZuS2y
yNIGmRFSszM+7y4Et6JJoKUhu1wB67abx9A3sSaqQkD2lSupCGG4pYqv6X7Js0qxZjGk+lB/5ER5
EwETva3VmpB4AA5B9UUkAmbU6d8BBt85EazyNrU2BUR0tZyolMnPx6otED9OJTjG5T9zPpSq1AD4
BA5MmrzcGapHXuJwKE1l+kQeFlFl+JBNcn2IICW35V6hYjxh1PK+6ysYXi59jUMNiGmJAnf+inlx
bbTBAjsVQkgL9Awf/jgyauin6IzWGmi44ahHURKhdqjrKjLAPQpn7u1XN0cI/SVaRmyxpInWwraH
4JmzwWAeFokwDXDWgpRCKk8DmID9mpzZcfgg+6yeDMmDsSGGOF/VwGLUURDwwTpLIFQwybCC6DGc
r0DPXNajrjWm8pW+FmhDKLsJlx7qIOqo28zxabIhtiIlXNKtduKw/+NlknTHxlpf9Q79PWZF44Z6
wtxOCSbVJKn8Cx2csApvjsLv4msOTPL9XHD+egVGNiFJ4wCc4DwS+kLk8xG/PEdPS4hKV06K5RUe
cXpYAh+4YHfpw/Npwf94J7xOYoIVKZIk3YPeRKwegEFheexM1ZnYUdBjfvDIGtzlovjIElX+nZJX
kYbpUj7aQtcVUKK3WyAwztXn3G1S25GSsr3vCEY/PzWFWgs5ww2RsyMS3goi5jowjrk3OdVUUn1L
wYiK2XiobYbVxrsgsKE4wVk8xHe5KpCfd/NY5zqV7nkUMEZXb8pPaEzNSyXhDyLfE8zid48Mn5Ro
wPG8gKP0PKb6OZbofl2+aP+VLa/Lu8gM4YALP1fY5opP+f3yz6EJ7DgRrnzI27ii2SIiUQEwG+Oo
7DWazmSMy05azeWVmsgxW7jRadQBRGCsRYmw+UHXbaYsrKfRyAQdQbzjiNaz72Whs+bmXgoSigA7
xozNGwzm8H09aymSNHtn0/eIPso006VSY39kKaFu9yUA1lq+UbAttLUzTTH52TfWUg/Z2XB5HfYb
FMQvij81m8DMnNA2a0/qeJuc35OZu3mUVPvz1Kcj/aoKPfttFCTTPfuDdxrNPFDcT+DlKyEb639h
LXXtUNOwLyGde5TZrk3QG1OLHICv+7HyX52LccpORFUE7tEWkhgvoJAEyHP4RKtbDUVpEfo8VvTT
BQtF375ynRuwyxGOD5o/Z7G9/mlDYb6PPccw6O/xNZQmRJQ+ebfyCl3qSyxev8ZiR64Tl7ioXXsq
JY7Cn+tVEya2JRylGEfQCjtPWT6y9imZObs6Iws8Xyp0kslCGRIcCHaOvJM7TfinOWExEYnOzsaL
qB6c3oQQDTSSkdsmAf0cjxkDZqgJFRSf9jV63Ac03uMwYwKKmR9ReuPhfaidNoGo0CP5iHDKH+uB
/EF1HapcwQEjuu0xWEVur1tazwaugreq+vWlT+Jn5cgVCSZ/kY9cRLr9pjfWBsu4UX0OenoTbtSr
MSJ+ZTEVZbdzofzh4kkIlzaZl4wVLqLvAwH66JpQqnDG7u2vHixtx10J2eg/+R3cPOhk4/Y/X67C
/bzr8AwqRYUPnC4XTxUmtp5u5GxJWPhqx03TsUYzb+ONNTCX1O+Z3jzYqXvurJk4e8dxPMDJB466
th2Rre546BHrDj/iT2kDRDNNbZMmUTEovGHejjGI2pKoPI1GUHFMcdiuGDMI8dhnetJd/xJ5Ck2r
yt224ZF0DkGMHhAtHA5zwGRrVMgTVhm/n2DHVaMLqs5MEQ4lfty+AwHDxYLEDImGRJSbY1kIEy78
qFVbbcmZhVwyySV88s3UGtRH8VcDiiwUzUBSFfyDGnr/p+tNIkVAUhavEvUY9C7zLt2AQurpEK8V
OAxzik4WUj0B2FHNtoEUlFz37wemKIYRlFa3Uoq7Ps6O44/3XLkALlBmeJCPQKvHEHCVODSiJT9i
hOtQmJ+6Nuow/1i+2hgxzFJpmc06c8dP/j0BbVzNnkANh/2NPKRw5qFLlCnunru5FNqlmLayDsJb
bx0O6QUiweZQ8uTuGrwIF+Jfvc7/LkwB7/Lo1JQ9Qkgkkw0OLAbx+HAS6SKVAVmG+BsOK6qmSltW
n7qSGHxZiAtfiBu+PvaJeFKkHG3eLU69SqrVfor4miMAV9aXvHHSDZQB3Ws+RyMeK6LhlDR7Hba5
AOIgfp8StpUz9M7uQUOA+9MS6MzzH/TY7FeS0XYXI9usmSSjQxYoL7IRcW8I7daLxxZrITFKpFAg
a+FTp+BzzHELvAItMZHQ5b/8nV8O+wdfYx18SSHcybgtv9PuDfdlteG4/iGuFkh9YXoeEnd6poZa
6ldiayqYIkfzFaNIU/p1YEsj/87wcLRcCvEQa3W+PE/AuGNwAjYkqEObuBbmgHIsMJN8BlsJAX14
YBVPAvgDNvh9IGFtHi6ehOiBNaQ3GAge1UUOJlDOR+18EPQK3ZxBeKkOFFyomrSVl2j7VtralqtZ
1HqxR2MlVdNUZ0Sdul1qmx8o0e1dfD6fbTQ4JG4LnSBlyuaYDEa51ueH4wO3V/7mtV6aa3y5OlPs
2GS+DW/gAGVFYc2PXQ+WkBAT6BJwDFKnOL15OTNGVVPCgnf7tJ+aW5wKabXiJ8iYhrysVDwAi/RD
siZhQbeo0INaUQcVizbFBec1XbmA9F7kUbCiy/MpZdkEVtGKElSxAgWTU9kr+7XoDeGCAUoABi5S
2Z9zVZ9aFTR9sCLo8ppO5AD68MWQ+nYD2usvm+7XwDRKqs1s+IpwDUBURm0dqmtMCwUKIZThdOBB
e8mRJbnxnjzZmzt23VZzH53UB6AQOouAO4f+RJKJMYe85vHlpyqBXvBnnULzeTQmPzw2sCNFZbJY
bbO8pzIxLZiO5oOtcgAF8RiUxpaKYBeGF+96HXDkb7oyQGlOK5SQa4JrRWweB3TEU0DfRFA4Mjyr
hvWNMw92syexMGEGgmt4xU1riClUyZLm0gyT1yTmXnL80lDa2hsUVwC2VITi85ZcgCILuL1iXtiw
MvQOJPgjOuJGOdspjUFHhlz/Z19KeFbtZYT1cclJPLtOfJR8MSypc5tJHSDRmo4Il0HHcS9DMY1S
qBGiz0904kfhsBKXObv33RQ+YFiusT1RwTl/nU6rbHpFhr8gW3XH4VnHCh6IxeP7i37MfZN4yqGe
t2BwmDR+8UnoCuO1wDYzLNYtUiSMLDRai5sr1CR1Qa9+RZekafA30xVP2Frl9tT/K+bw0CU9cMqj
/8ZYEq5dZ3Lr55vNbcx7EK2ghVY7Dc1JkX5NztBHIFaLqpWrwXvwbGFgD94MCo+vV2P0NzkqkRiX
JgExTk0ys78e6CgWtbaksQS60jGi8ctpV1mVcMqBz6TQ904k4OAZb0hHrgOug6zh82IV9sb8DIuE
7J1MgwapyzDcnA4kNA+gUz9WmzXaEQLj3kbNIull3HA6OSC3PGiVgMcYrBnC9LFUjRWBDJBvB7xg
CxE1+z5kTV/AWuNVh/8Y4nhj5QwUzPo8fb3TtpEt/rGRHE/lT2Lyklzo+5uO84+38Gt81g3m5Og5
gWFXR9uv8u7bZ2wWumyn2r4DaoRUTeQfJDp4pmBF7qFuP2s5Gaw6Bq6oGhD5U7y+w7paXbL5v9vu
m/+D0CpGLF6GoBHJE6SmhSfLzewmNalc8H9HS9lwa7LTA9ORKYNyOm3AT1ksy0LQd/J0wJFbplKf
RH/0zdYv6Rs+lDphGCnO9DuDQqjSIcDxjuClO16DquWbXyydGwutliPqi+zFD8QUOqAVhbUprYjK
/z/aHgzI/nVvV4W4O63W7dQCzehJt+CKoAI5TaD/yc4wCtgy9BST4Omd+DC7OpdbFcQckpwy+Yls
IJ3PbN4zlw8juEVEx4Pj/YEqEZtOg77X+fZMhxX7OAT4HNrLFKlkxPqaq3DLIuF1HaoIOAY6eDF8
pf9kcRMPdGHauMv0o5SkcTE/tt1zXVb3OsPheyiCaefskLLy4sVWjR89db5e8P4SfzulR+/pGSst
o3+1+Dl6S35NCU0FepCnyd8wqOD5B7YlcYYi67NqqaoXE86k4vX//Plyldu0tkp6zH1og+TpyQXR
djICQKkZEKIMNJeALufo65SOcB7tEBqXxYMB3P8o8MLhIApxxYH10oAVu8O7Sp98mYvH1YuI+Y28
APiOWfHNQTeJxJYofmqLFey5EHE7VcruwVeKQHb2TmFi1lO4umrtJPuV83Bzw2ZXAkB5V6thQxrJ
oKnoBai8b0Kyw1vlF9ajzOQG1OFoStiuL0I27R0EbHqvkPjZBa3bJM+UMbDnHqahvCa5EHUEyPky
KxRWjbRErBAz3WnKX5KhL8+77rtfgzpNosVZbjsoXP0pHVBpYyJ/d+7q2jjmEoVBlzzrvS28sdDO
7WIks6z4CDzAsqUWptpIYYLiYVgFSf4IM5oVPWn1wNVF4VeaU62W2hyEiTfWi6+9gFQuavetHykr
A8RaEMhOLocQXj1NAXNI3Rh1uLnDYz0nzE58P7ZZNGLQ7QU9ilmJsIZWG7+lUAPDeuMEkk5eFO/Z
3tI7MdSim4IvhyxdG8zq7geBzfDBuOTnhH98MwMazWxIH7lsn5XYlseoji+aJkFjTr7SdI489wdu
Tm/+304Fg9HfcGkvOHjVXKvValvOKTgXMKSO9ZM1su2JCVY7486YdxlVyGTywFibi21qUmXxL6u2
u61BeK01W6l1hK47LpnOmJPLOUXu+r4pJ4kdPBKGwW/p0WuwPs1UZXwEF0l16zIHjV2YdqMiajER
uHosEv+bqbtTOW1SrA95Gqx5VjEnd2O+AxM7SYjr+0hIpgoDHpU0J0t/0WEWs1c9mac2InxJwtHg
d8/VrFtGmFU1U1l65WABFxD/0hNckVVNVLtf6sYe9g9ftAeIfkZdctlmupGpYKW1zbwrFTidNVem
Lckx0emU7xv815H5kU8MiveyFLNlUDDqrtKnvX7Is/dFhvKKY56KsgUTgrZI9f2/HT/qRIj2+LDi
fc41/dhZaxukZCYdqtfNkaCcL7gomE+1LAe43V6aa8F7Yve0SPNjm3811mB4Q3hgBijeVgA49Uz0
ZnQBmEIhMmKpuQqg8U8qPoCy0/py8dMj7jReawjW4vsmtRZ2inr9BLGNJQic4P7JuFslSPcfYGYn
q2kMzYptPkNDxZrYy/D8T/VSOQD6/ERHGqVwjujXypm6GEbBQpM+UsqraDmHOB8Rjjqp3baC2Tc1
hg0Xt8S4v9+siGecOl3ilhxUAzDsolk2/hW07xIfYnfyVup1dZZgKvP7kNMFLZxWi1Ts7acLXky0
GLE0GLyfBe436YpCGZEFDt8lzccRGJA0gAYXZrcZo9X0KtxcAv5gku9RPaqAb5YYwHfC2KKU9mAq
pWNtfzKiZkwfnpbRG+WlDh77805t58aUZ4wkQnifvkYRk7Z8Ju7QCQXY7nUDANJWXwwa2gXsB37B
PkK6aAC00WKefRTDzBJHCuITCbxfJh0itK5LI8mezuTB8bL/CyFyZiFk/jQxH3xpiRHwM1QcDEtQ
hG/xvvQbJ7ppzxIRr1djrxeaKUIHjnFn7ItdxnX5Fq4/uNWlG3ybUZ4SjGwuz0pHFsN7kVn546dn
PMG29cIFvWNfQzrhdLWF3IzignK0d3gcN65VpuQgbv0cdK7/BCE1OYCiZEAP99F1e4zi1KPzivzB
vhOIS3rE/hA1aesosBNPMTfdnVflwYnfBz98AJYusamOJnyh0SOIg3p3VMq57BhnLvqQVqIH/x0s
OGo/vpwSHxPjCbjmS/Z2gp0lSzlacswspU2v0DcC3FuhsFQxb36YTqUR5eYjr8QBUct5qJgSYgvF
66i1v1YwUyYTx8c9WGDtdH5iJawEfWI5LTayCoSsViKfL2ZgQy4qw1Z1GgKFxTd/CN7yaAJdd2fM
riBudIf8LIoIJWUk4LWpJRE4T0ufEnNwngOwpp9f/LWJjOfCHbZsbrFCPoHxjTyYzbT2ON6jbKou
7qG3IXfX+eOpGgLb9FW92FozPR9+V5NF7InBc779E5psuxdXvdyXN2J5v6//K6ZKHW4FEiAelras
ufHzZu5YW4D62EbZOOTjll4zzwn/swwzG2QkebHMuKgZdKrfPn9PwdZJgIexkz7ORGMrP+2vUDKU
aKVWyjDgL3WFkLT3UPnY0NPVAXPMkRjoVVnfMDJovhTpRWpnbWATNWWKv3VeOTE5x9HHEmmwxdIB
eZ7poSf8bnXC8xAbo3UhX5LV5JZgtQUI7b/WJmGBNzKqyJVCx3uBwfQdaWPtRmRMART7/NUssECh
5+T/txWoWQmc/RLxcM4gVRE6e8D5O5F8Ah+dylJuS3PnIDWxFHozN20WxqyZgea2S+6VZZ8lvtvj
UpLwEeqlYAqHB8zc9uwFQFYHAEwPkyP4NpntftYbOjZslj97mQ6nOn5ggWICummy+ezJwbW82BDa
1qJ0kubpd8Ka66WVFz6MuUDbZMhUqalBYD7xfUVWIrEbuJ0aaOkb0eM9jJqR5rW+Th7HcckHBNBR
brHscOUX/ky6zdbN8Jn6okpcp1jHU/8PrA137aK6L4VxjvZGZTTTFWiZyOm1t3l+9NqB/eQYiFuq
1pXw7oYCICSLm82akaSiDCvfVWS5mnfQlBDXHTxy3vFIBo6GD1W/szOqPK1pjFBq3ahXYSe4WIa7
B2x4XFIkK3iWGHWGSDBoDvN99v3XOzEPLAfZ661HylMr8VMCEwrRcWvalq6X/QIjC/4ZIRig31Dv
lRiJMStQ07Kdq/G3rjjUTmsuxbUaz0ABkghJ2hzozvXnXnpc1gQdxQZ+upRAQtxj9/l6iWl5+xgL
GPLYmlZjJZt4SADqg17wHga0fqKhwztC0wsh8pnIwumh/4wbbTCn1RrYX7boDxd8AueK+GSNrq4f
bGUx4LvDYOMH0ZAwCZV8WI+p0RuvGgOOFlk6hVzx1iFl/nK3K6BCkTh324nbvY0JdGyY0JCj4E0b
jHlxX1AuyUOaKtLpsChGrpSiNu87vKjefAJ90KhUh1fdvedsWxuU3HjSI9oMApNzJRYxVWCslmL/
b4V8z6QLcq12nVZkj2zbR6iGbwELn3t37ubMZ/7ANjunRIekb/a6FBLdZ/GrmEPgZujlcI0Jx0Cz
jPvPwETIoCv6v/BGSgGf4fX7yJvFOMoog/G5pc2P1eSxZfr/4epR9L6txscRDzWdFnVaImF6nn0K
CalCUSe1s7NBhKypWyPnh82CWO5u1rrWgkZI6krnZfLTuxDuF1Ytmo5MwR8mdnXO8LmzVMVs8pX7
rXy00EzylYg9NGwAhzrJgpKJKm7yOFGVoZouIZBjCWONOZ08r1F/dzy8EW/JLbw5BSVPYyZP803u
sKdyDOr21ROHv9mi0M9+vDL9J2YX9FqLJUtnbqwUX2eGWsRcoNQPPBb7V6L4lS8eDuu4TCd5lNYA
Sdr8G59NjgKTe0WfJFPR0C+tydDbqXThZ4wms9ZcTyaQttdaH+r5qd0ZdNdLpA704BsiauDTxbpX
GebmYKooRUtj/EQ4Hc0sqt4MZjCEDYHA7Pw5j8/1+2xAYjQRgrjYFWm6YioS0+3GTqOlhJhNEV6P
pJzsQKxtgLasK6KN8QQ9ykWxXMlVW7rNJsN2lUPMpuj4W4wsUXqAZqUxgfESFNPJcuXo91hOPk+f
/Z16VV8dP6eC6qj9eAvvpjL3f8+tHcgalRjC6gyzRC+hiS/FlLDeyY6tRk+9q7hSP5pVIjmH2gB9
ghvVOjrctF5i7Ng5NW1JvGzvcYsDUWIquMC5fo1ePjkXE7Vuti+90185fQ9IC5n4st+KwvM+kUJV
BtIOjt8tGC1b6bMG4eoQbmgKnHHI19pOCrUnG2NEFLv0oBTEo54I//i7H/1oYreTbkyNuaAh9j/z
LU0l8EB0KmGmW+CW4f+l5UMdxlDwo9/jlpAyB2iQdHRN5eX//ymeLX65pypFrlDYFwiNgF5YVP+8
d4M1I5BO8UVUdThdTn/U14NdwxSG48kiu197K1cRKUum+JYBJu/d1iRkTFuZOEDx4alRZN4tqSmc
lMWKTLfGqfhMt0N6c3C/MX6pZiwYDcyf+WwHuOIDXNy1CdLRRU/tljXmsA5AeaFwaE4cDaZux3NT
9C8AsfGI2AX7FrDmYX7xtoSNHbG8HG8AmlDt9sP6WR/zhTX6NeGZC2WpNqcphdtGkxwYwbmrW5YT
C0qB4n034vcUVcgs1rDJPy4tRi3mzdeN4IPBX/2fS/gmfZOpfTniOpKENAQ4MEsKjLbvhaxDZbt1
Il8w7QXN67gAeXu3ed8vg6Q7uhqWgt/gboJHMkt6wEE8d7So2JQrriUQ3KLFevK41yleH8TGEXAB
9Z5zv1NKCfpTsNu/402Mc7+NDoUjYnnFnQMLcU6NO8gI4GPPAD5/ylbPiNvZxnuDiilV6wxfOQLn
0OyncO1S6uN4Aw/pb8iJ20CNHeGqfmsblSeQbbMTN0/eCcOMzcGMQufRZ26hO5D2l1MXH5JaomBh
ksaKTPZPv89fRA9Iyy5mGTEIffI63d2dNSYAzk/Rp2MlEAnHJoG0P4lLH6JJ6cXKROZb3ixseROF
tOtzzSHErBqsW4IN6WFnjfyzB/gZqfAq5V9wgqmRt2rLLZhMjLIeZcuJ/K4Wlf0xvY9R7KGkiAc6
aZ9s3BGmDBY0k/ypJr1nL7/ZnBX2ynAe3en0GBC2BUIv1FtYH9cVjj5gkDCrfQxDryUYEkhTPY2V
ZX3PX8rmj717GreXiwcfLZkk589F0rUzUh9rZw1a+eyXwAENJSaBWiBOKuEKoEswYwK4uQUBDNMc
+DQptW5/0cYQfLmEdtZPmnixfYZ6ku8Fb3DKckuYhDqgT2x8K7+ub+4ZBIRb6pIHFrEkHMitrQvQ
sXaVsMQUPF95Gm8zXAcJ82pJWpSxVuPQkGi6imgsR2PijmiGhBrmUIvR5jx5uO2H2S5LjaBnFO1J
U9nGU+u3ZtrPVz16vjY08dhJZBJwtpfr6mYUCEbHO3+WXYdNd9JkHamsQd9KCctAM+4+6Df7WfB3
mSxdyOzT0orEfkvTia4kYxzhNv6g+iG/Zu7AQQQeRUX3Z3zugdCb7hGr1NI6tXzaGoQRz3PGaXp7
lkwYM+LfWaQF8oeJI8pcdgDaBc2MtvfzM4uR36wtPC0pLkiMdxuYoIOL3UnDsLaOad9VMxokcUrl
xpq3U/krtT4dpBWvd0NBgOlaFTawbLSoDnwwq8PuFgQCprqmbp0y4OMrbo6n1HMQCX4FcsIbVZUB
nGAscmCau0AJ4JHKuqTd6Cvhfybsd345xCs+5NOLqlZkoB91gAkqFLYp7JtURHYI4Jf6GymMzUd+
t9XIlidlATRx9kV0uA/BL3p+Ynd5AR2/LdxDveSeUh94sMZ4zR+ChGv+l3MDMSJcMUgG5LGZva0G
X/qCl51/n+w6CoeXF7CSwDbgJ561T/hMOfzi+qvk/KseNOUWsacFR/mseeLVfyovGKjuJO3IDAej
G+7P02lCC0pnyNTWE7K+/2miRREvl0Q+sDlchngpf7HmLDkvXLDsMJ0lLFRgR64eay2GCYnXqkYN
9563piA4a6MLghV0bQUZzLWQPC9Lcas7J2iIshSmLeDmWulbBTAPGo7fcOukQ9dR+jsmwqStFA0m
b4JcHrDx0dh3ajWXSHF/uh9dhSzEtwpoQuAZJbKr6ppyeu2ouMvOqhSOhHhO1Qm/rX2jcop162u+
NkCh2j9fNlLel0Ud38VeQ5fsq5SPIvkRIQua8ebnIbZf6bGRhXhuKfuaD78f3vRMF0hWpkt01tWx
Zn8YoAVKY0A4E+FmusoF6amxL1ldK1zdvV9rRpfudD4t+/1eazhK2HhUxxS+ZF8gy1YW95ARzrp3
04PrWME0iC5SFfiQCfZahxoOXWuDJvmLaq8V+ApCIQR8j/SwkcY3S98cQOAxYyGWONYqYtlnY7Sl
5VZVlaSp87YjLGoyp/lS8rVZprc+xVhwXxM6kI8HMMNoTKMXVursU7OAykZIHqF4PofKWd4lePOo
mB72m9fwhQnsScjtpui2PWZ0M2MBJu41gYZ0/VZnhmNqO3E+i15Ru/CXOqOW+Ua14fJHuViUiEWb
wxmQy9FQR1bcKfTHfeykhLI5ZA+nCf9GVulZywhLHRNGRrBqu8v1xv8+VxeXaZxyawA8RwO5kTDZ
ZKiYxnydHJ3HeynQD5GBh7RaE5zkVwi14rEhErG/6U21JUPtRiwmWe9778MKg8owflrHOwmGwgnX
N5pWmJKkOnAHHJGn+R5jzPcASdKW2dQdeiTnkYq2l5CPJngVn5bl3MptHw54Fz3jD0zWBXUIZ9HG
QCdW7VOUgF+q99bNWOjx3NgLFqQMHuWhVXwrFWipJgOalHk4c5FkhryoiYYk7T0Zin1+T9bTKc/B
6T5DSTmNWYGWutdrrRZExNdTh7HUZNjFzhpXEakrO35RZel2fa7w3l5F/Jjc5oXZw4MRJ/gaKkm3
ZIFvB17rXGXcy5YSPrhbndAPate8KLa7NXf/RiBeTJaahP14TX49UL+ldrgR1j8+3qrQzgPA3vZ0
m88ybtyofKc5O3n2szebRorcMz9S+9D/rxEAGmOUQhj3BECs+/GUufl5RStS43cVXxsrPLLdkY6E
yvoGWccF1Y1rifFLfqfPRhsAY+evWDRfmyi364wF4XYagJEdF+41UrTBNjDsIi6ee3/NpwEb4TfD
KXPY9yH5Tyzc7rNPDtCM0psimVLwZl7Chdv4uKgGlkEXBIa5EMgpf2QLnlZ4toGhd7MVCOwuNa/7
G1LtkHqRzMn6TxZQkzHFSx9+dDanhVvvToeOInbxK5jZaTm3hw//2PkfudTlSXu+4Nzncdb11ggy
73ulF1z2jJ7O6keFkPEY5QRh5nbJ1fmBsVfh4DeRYO04+CDUBI/jsWyNwyDGFYGkN5l3LiwuiNgD
47Ib48bkQHgqXtGo+tUgmtHYamYbXmuJGU74gi09jfVErJHjxxTg3nTUl+i2sYLhQ3uJu5LPKJZA
NkM6cF+VpNa9oEN554oB8FCwxxDEUyNlQ9+nEDuv+MIXyPUtOsEkdKgLB6RMKU35edo3sW3zU/Fx
sZTi9jXUuGG0qCHhD8FYnyCGkgpUbDbBvZIbPdrMW3iLlXDXAnUUxgaPk1A/WGACIMyIz6Efod87
Wn/AW7FivGjX2KQvENUy3I5lHndRP+BubOOzNF9Sew3H9Qk1Qs/bAnmmAUCgxh4vBaeei1JxI8IR
Q6d1vLUnczibHFa9vVWfwczjBBoxYsc05PbaioBoBGQ75GG7wRT0mle39PQKH1s+zYRAzZhKn/Kr
rtireKgNyJJB5NKXYjzNXWvh+aUo/wVkKoa1A85fdTuAfNr2d3dszRNvA0HNC2dcfAwH3RjUxGr6
pC/oea9jC9qHwQIaNDjIzuBKifPkEm2fZafsOUKZKuJgQ5M8aQQnehYD27T8Td5++l+EvsA6pU/v
z+1bi5PCmIRYmXnRBHNVBsyCqhmuzL6DTUWQJVLO9yjBGNp6RI406A4N0WG1bkbOe1w4HeDdDcYK
kCy82QNfW8grYACPqnZcw6Ky815gWX1oPRhCD2txXYGwiX0PPq8W3V2qKAJXx15gmzPRIHnf7kpg
O5MSRu4LTa1FQ/ZZr8saIQRvHTAPJnI7qgDeMnZ3msD8hvkyAvVegdBBkw2aQ+HpO58YOqq0X7km
EtdnAEe+GNbktK33TkfW/mW67PikRW4XVdg14P/DG1N5q3OTV/Lf3f5G3sTEVdG5qJLwGWpmBAx5
8jYAhyzgvsqCZOO+MT59TkJsquAW0RKwNtwCDWH+FxvVFlB+tjTULz0Kbmye51FIYHYqhmctDmVZ
Fadyja/Zr7f0AnFU9rQHnjJ9sUpZK8mu/e88AOm2zKF6LqMPMnfhLlDVyBHLIztlkmh1Es2ze26I
uDcUSmxFWAm/FMU5kPJgFbf9wR5O8Xcd9iiFyphFWyr1o7oXJQT1nN7LY53aaED8sPYPqpEjLzr7
aDJKK3MtjRRGtm/pWcm/2Huv6IwHHAOay/4ShwwjSCS1sFzKisw9tb0xAgEpoufpDItO7FOO3lM7
cXNUMWztqVqs2aa7UBVz+yLJHudFTSAWvmNO2hAIMpfV8qvV9bqhd/MzuOvxZQ0IsV5JQn2OfR9Y
tMeXMlyuFCqF3aiDGfT6EqC6Nz3JSBkBDGEF+rmbHCeUDb8A+98aiiOOfplW+cLv/OwAHupH1Dt4
lKRvFZV8RWmee8HESrJrIz9PhZGCGYJVw0pIj0tSjit76ITxDXDM2Pc2TrRbkA4FVMk0oLfc4NzS
tzf9XmKUmmlHo6GkoVgqLmWI7nE9+HhkRFE59+au3xXPHUg7dpdJPWjeEpwApiO8lsTUfbleu6v2
x0mG5Ev3Sdt3jxGDAsYftKwI5IN6y4OK2kouq1qLU9Nhj7rYgAIBOj3zYqypvWYcPyew1OcMAOjB
vsZjlFYMCKMkhaiAVOqRgjKYzWYAHaluSUacUj7qhjQIibGkPVY93nj8LU3wXfkeMY51aLEi4XQg
Tf0tzW1S2Z886AoOKyKEV9VsmUYM4AQF0jEx8hFaF1d+eEm/KZaVEu3rmBk30klwiGZ8MbK3yVna
pWBcRv5RKvOU6e6n08uUjTdcpEF7h95Nz+S78oqSb2tFvqeR9lRYRqAWhy73mfh7pcFX+QvvSG0g
xvQBJrgTI0H3ppzqgSHaymyuhKgr7Y1wwgm20NPTTGg4YcIapHY/HDJjTVbBaVT0710Vmu31ouyH
w6hWTzOE8gYuHfFnq6proGYYE5jLchHA8OHqxRsIM19jVE7yK60UqNN2yGQ2mehIXAxwxkfRQlBN
fU9vx/CRWMPxA0yZrSbkJGKTmoNg70FBl8KgcVt6qYuT8jTfL9BH4jfT+IoDGHsuFLXaEuNpTnVT
3/H1VDsxP31BRda5jtHXSK+LNHKfoGYj6pqSThQ5VXluP4wtSNdhWYLUOirnyjvulI4aQKQAmuO8
eNJo7jL2ckyqEj/uq2gJAF7jRkXaR3LDNk2iHcNMebNP9h5QCqKKjXQSxmwtaqV36le1re2fWCzO
++TqCD7eduo5OhVYc0GXOU+ORTgO0/Ci9FPpcM/o8wy7CqSRDgkP7KDkJnp/2hJHdht4XpK65aFR
gzxSwhzZj1fmBJzilZdDUMt0OvZb5LEAMCOlzJWqVPXZKimvNNtxseUoTctNkjgg9Uhg5G4dF/gj
gpwrodpYCcsNU7U9zUtqoFbLAUmUHr7dnXyw4rM9w+MnHuy8n77bexM6yJW5DRaTB7cO4Ll8prHZ
f68nxg7qLhU5qBbyxaY/aAIdvXnvbZdoCvnYdbk75V1NRJ3ig/rYgiGUxeL9vtbnW7KcJq6539rJ
uCb+LV+3s0LmMChuO/IqggWIu9n008bs7IjEzchJzpHNFZAneLrmyyH4qUHY7MGF1RJPfRBpbtx1
XhkWVzSP0cMdS660jcXoh3n7IvsXOl9yj5a5vOtZyEKcGpKV/PZWKclug5xcHfmJHJqQLBc846pt
Ir8QuH4C81X0MIQErHkeQStt7whCgYe1rxLDCAi7KSVFr6vRwU3C+e67EVlmy4NTTQDEOvAU5d46
u22hHTPYoacSZzSzq9ulmXW5GIFb/A215rW51jw6TxZMQ5Uw/3DG0cRZeoXiD1k0lq2BmXNIn/BU
BmbpHWRsnQCwxiDeKfScGZV5jhkYvOoEBAmn5AOWzM4adOBgRd2SYlyrDWCkKJtwMwz2QlMpSqWR
1kBd1HBUJjtx+5ON0SXOKNXmT9a9l8+2IcXaePts8jGhE2DminmGbvKwQHQcuH7Jx0FjlMgGz7Ww
Imz3eLM9NNSh6s8GwJBs5JKr199sMtYSCKnLt2Ftd+bTVYZgIQz//0tJCfZ7vLb1Bs4HGfS2p8KZ
zCbXp/GlcA4cXqNa9yjFVn9YSN/S6XEB77XRac7iqfiPZSRByz3sbILTp8NWmsgjBkgC2B52mKW2
nxiq+Rq0U1dUvOfQPm3+ZXjXVs+IUWIlqFHXolfxaE1iWiGU0kCtnSn27tiz6tX60V0Pfj0BzfPl
l9IrmHxROrO1mZrNpcEH07cDZOAVVHulXhok68JP0bP58fyLXsqNaLLwRexQz0dv+hDUp9MxBXfU
g/ClYAKwLLfICxpQtJ4jrzohRBwaYW01FjSP3S0w65Y3xYAqAEWOgg8oNYIc06DFDyNkURFNaJ0+
dkdP0zc3+2sA8lsig46anD6QgGJOaWSMN1dHIoVVS5dGLiU/h1eUsuAZij3vecrAXolRU6CfF5Z8
oKg7am2C8aqxKgdol1+e+4IcflZNC4O699XiZUUGjrUuInk+3xoK8nCR9sa/XMOFQ/e9SRCIQO4a
krjevHQ1Wpfn4QMpDpZHwlbTn2EIADjlnSMh4M0KHXHJHKPphZpZSJBuFPa9SOJimKhX67TPHguT
bICVTpe4YLqRKah4ECLVCOctCLjp4y+VjlqMyVkL4il5IyW8c3ltbMUgpjCLjuUtmTbiEZ0ffD+x
WG8gf6UOJTexMELdQxgRHhoY+tgFlfeqzAGG9Qv15EnpYwm3qEGiDCehUlKxH2uh7jNr/Jrkpz35
bngNUJkYeHObaljD/Nk1L46h95Rj+UcUHOVUDskvbhW0Kxz+GZ+wcPWlfev26ot3Aa67HveW9ei9
ppqnOkv2yl8YuVM11q/wTzqjZS91eHmVwkol4dRgAnvd7y2P+0VqdJ1w8rS2/BOwKGzjeS11DScN
ad6LVv7FjLPyDqseKSbHZcEjOONItppNUawaXBXOFaqUQNac7Pp0gCVv9xMorkfkXtGrpZFR/6Hi
ZPbQrw8V0ALD9tYmfJdp7ZXCatphkXNNSZWDkGaJ2OoBQmmh/mS/fRhaPPnkyRb6u8XTEzvpBrBk
QtBLCsCi6xAIu/IZKNUlJQn8qF6RIYfuj7wfDDOCfThbMxT4q8GYrZ5ex/1uHdrMbG1amrgTc6cV
5lN/bC0FKRKOP8YK7wUihUcTc41+ZE6FybsvY+hpYrcod6XRPlVhTKlAcE3oWQKFsysrlBrb32my
5JFHc/Sj45b4b0llAG609+M3/2oBjMOuC0St22c6YQ48Vrfv6xfxxHaHrTppn/yZ8iBfdRxooCUd
yP/wOB4DajISVC9OgNxbYPsujx24F39gOeB2sBbmQCbLZeXOIz9pg3Nv1hR6dma6PxMCgJi5rUIJ
0CCt9ZtNEAAnv38bDZ3FZohGrzPBBrxfn5ee6FZ3OyoKzMCvr5uxxo9aVW+6SDSqzU5k7ChidqdI
qJYJ1KuLE6DEZ5+9dWEZTWsnG6cToXQ2HztVFIopjrbpBu9cGvR1ano74DUf+4CrRJknEcHg1ibe
Y1JQ+p4TH65QuZM09PVfPvVhETFpMHFJexSWYJKNdqd+5l+7dAFkrYqAENqqOu3Bq5EXbjyPZWMz
VJXNqsVC1FylwZb8bo8epPAd8uGtlYeVeD4KQ8saAJedQCI8kun0k03ca37qYaKdMef+LHDYlE36
4pUX2DPI4XDFEBV+SlRymVeqOrGuJqr1vSmWAnADffK9yzzYakuyNK11aB5gszt0oGPelxZw5D7O
KOwWft0WJn1Wpb54GG5UKp8rvibO6PKnX0S2Iri9beSzWJLmjymtH0pWpnzDSxqnoAVNAEYteEAC
+tURZQW3JRk3/iS7OAURgmhPWzaQIOiJn8sJU/u7tUd7rLhc0eQRV7RZmyTvgYUeHBFI0QCnbpxQ
hNkO9zPwLcZP43rJf9mGIl8u9xQYZbamnwToxTI2xRUomgCh5bkbZpYoLdDOCDpbAOdvLXTu6la9
Jc9tussd88AbbFLBNjZnNiU1yrEs4yNc1n9EAX6GHtx4zhCvjCMr51JGVlamPmWRaj7LViuDsjk3
CwdZWP1P7D57/vcNOTmy3xpzlad8DFXIek51ECOXoLq/N4fhScHgts1Y1fClrF7aLTlJ/kpvvRQw
qhMzjeFWDurbfZvgdvRWxv8NT4JBNrPfpanYPWxBx20RJC5SpxqRzMqnQxcHy6/edNAGjJGZAVXS
2DqHcXjcKyD9VCN2+PNi8tXMGaxyjm76Kg5wvP8YyTKxpk2fzWOkAaZxuMX5+xc4fHk9M1RDa5fY
qUfEUvXg+swk2wmGil/LiJ3kOD9AbsDAFa17sfp7sBIROP5j3k8VRVIhz8pwc1KrYn/HTSyelqwG
+0v01rEuhQs0K3OBLNTfnFKIiHwSrTC8+9vWju4t+SCF41LZ6I+WAAOZ5QrlRUo5WtwL/euJi7eH
jxfgr1tHVbpjT087oU8GzNzrska+J5/O7vLIDxZUAbnc8TOhDBRXlASwI8RdjSXO0SUXfpcmS0zv
NrhmTTfhshbVHGk8LtSPISxiFv81sSqrb5QtieKxydk1Dhd9GmwD61Zs/JkdQP6U56RdXT3V98KQ
br4Q0phmYgFlr05dC9G8hxVmFuimhKsX9yMfELc7f2Pz5OrQMwo8B/TLzIHvVpdz6Jd0/rDPzvCE
kIi7YalnNo+5v3YoXtaobTdEMqLXEX+VlTgtWDxT2/f/gfVFqFbpBy1W64Jb8SzbnsArSv8xZ1XS
9jpLJVRT+qDGMRWpkELzhx4JAU5KHI3xTpP9ciOkYCj7nCF3pbRtEkReYrkhhubp9T7319DUc6tp
qG1GXv38PamSG+ylpm0dK/rWPg5YqAgn1CA4AKfphzdPDwrT6sqcNTe/8QvqjMqI86N/ZUBRDj1/
/VFoqDdYv/hxLzSe72H5ueCKC667pG9ZgWVZksDx3r1z8MYec77uctuNiIml2TSPjJZAwrpZ3Qa7
iBRxZW1Rh43Zc8fko5rp2CpSGFKVf1h2sxYFv3ClV/DouOjYklK0+KFFjDMOrNpOfX9fmi/JLP9m
y+Z0q105LPnjd8eqjCEwkOsUevyWY5eX9vTbNfERlpn8j6B2KtGC2k8E0THV2SuF8f0fIrMOKFpu
zsuvVzIpn0KEzuPRmc6zu33fnVYhtLAkMzL10Tb4B45Offslee0Cx+Ov/M5CVyg2RHzcpHFft/wc
+sMC3229qbjoUvzwv/4wdymely5OB1kBV9LGuUQf9xxoet/jsl0qjwNVzlO3YD9Szl71CMNEDdGw
P23thsPyGvYUrSVnMNuDAv/kW3OCpVwSJ1l++v/DzZKmR1jDPwTV026IT5jzSnq+58sz2AiBAxhq
U/8NYMC+4RT0hgo1r57cn2hmy7GcBqzBrJMKx0uYyOSrxZ/zBvFIs1KznCKj7sUd0guHdQhqUAQL
iw25zRWKQ+vbcscLiVF2rGHuYeRKr63ZRzw7+4x0++/gQ4R9/EdVpvobsNdyu9wszXAhf/Tp2M30
MlvcmgtqPkM+O9xV+D4ZhhnxgDjnVTk+9HjpTQ2k4XABx0Rerb+Z5FZZxYEnhO6AJRwhMxINOIML
jlTmGQ0T85gph4uoeuSOHnpHrJpB0/oB508B1dq4UxOOa0W8JUnLjMFpccrAAQvSN318AZw34hTT
GE0RyAn1bmqu4+LY3kdAdwtKzS2GcANHZxhQ+viOB8SfRlBdja7vP4ulGeFuB+vlyY4j4LMz2YXR
8EHVYPqSV+TAbOm8kvwEhoxehc+a3wiJaChSOGVNuaioKcpqhCOb34s8IgidzayU/v65qCVyQERF
Fp9LDGxtlDnLdRhIrADl9rDZ3pNhOoEojhF/xxffhpowbkGiVDyD/pYuunUPd9QBkWa9tOTaTWC8
O7jZRS2JFkt2QEehsQbzeQKFvHhUMReUPXZWQS5TRTVlXuf4bSvaTxFH6RNBMxaFcQdA7uMfpAbp
dm8yiFZ3I5mwv7VVvC47Kf6NPpjX/2GtVOS4tcPMmthkDE8G9k7TgEhdp6c5fwgtBDMb+wC0GUBR
Nyzo31tSWt+V0Et17KASfCBRcriYb8unncOajb1cX2oXlzzA59fytod70L8GpnFBAKvcX1nTA5SJ
Dh7rkdDirPMlGAWAWlyS/ak3pFLrPY01yzdUI2awbw1stMWCv5jzANgBrbeibrT1vZifWGNyOyuu
LZaffpXxZpq+RvnQs8jya9wPNFULfzcL7npC5Y9L83XSqWeGOGOzk+XmCLTlwFpThzyeCiesQZDe
d8AJIx25kE3s16XyHD2JfAtzlsYEAQoySwdWLHgjwChBbxQQk1DlQDajnPoj8VcKxBjE1EJc/Mxa
YlBgjYjVIumHthDWxS4mECYkAG+rWE4D1xHxKfasswBNXzNNpeUaLaRovhszys/OdImjPuerY5ny
XNFCnLBJ0PZ5V44b69nvLXppYd45Uv2eDagvc4cQrq/kce/KhI1q+ZWm2Vpa1ITQfL9knZdXk6T4
v9zt8+bauZdquQeQhott570w4JQ3qiU1osiFoeclNMKRDjhHc3ba/KQbCeHyhiOyXoAbHWjD4dCA
jdiKJPAuOCqRAv43X6Ui163HM/CFUYv5CwZnYU0t3xJ8vjL8bArln5LdiCt/zw7KoLwLiC7O01VI
t5FqEp42NO1p0f3TGaPq2dWUaoTQSCZagOFekJAuszEPmHUTppx/RUpCFFf6MdLtvTptMKY7gefZ
Nxmg+YuAekWNgJWwXdc1ASxzzjsINTtU+Zyngg+hLfewVm+OSha0jLK77ePN+9m0WRhn0zA8Eixg
tmwl8JFWAo8jBVD42EqKNfELnD35+YNd4gklVdBd/LeBNOHFp0bn1+fbF1/4OpUOTSCKg5dAEm0g
NxSwsHwepihlezkgzbNcqQK72MqzR41a63leUxkgrYtK5UZkrDg5JBwas7ueXCYybeH8UJDFGVjr
VTevP5voD3vInBTq4CJajpHnY4rVU6JKqaosSWiQ8Wc/UWGHYqT9hATCXZYZBRC2sF5fD7fLz2MS
rF5Rit6YxpiWC8sSAN/EWGoCJy+iwcqh0zLN8B0ult9C536HOAhROzpDywVN5A0Xr/OPfziFGDC3
Z+LoiIHDvIrJhBgrzpmcFq4wDAE0V+0YbPXgU9iag0tsB5n0M9NKAGkOJ28ZytlrOWI4Naciq8+n
WkPiEfAipEJxcT8ReZ9QuRx07ZYf855zEEfNFnP3Jnihrgnf3L1pa3X7BC2cuWnA0vwg4+oFDp0b
azJ9wuhAaRvuDauO63UNbHIyIQlu1KtZdToyMKBEpQldfqdUoRK4+WYWvZIXAqkaU5nDeyryvbai
h+tg39dTZo1D7Xuo428+A75gGl776uLXxF8em21lZhHnbazVxkJ+d16cirPCVcgBoKlZdHEEXtJE
xpLd5Yl1QpLmyF/Mg+MGV11dvOgmT+VxMnzy5oDXTKPJZUJV1qKA/59eCSSMiJ3tgg/CvWqM4My8
hMKnEWpErN5z1P8ojYosfoqaW1IREzJOpd8Xl50Zz2ZJmoTDb3zXDtjo23jL37o9og1rSO0fhcP+
dIEjQqVFP1gR9UBGYQDKKduuaPIF70vcI3HyGam/zqFBOntmY/HYbECc94P6tnn2vZwrUmUBxfv+
5ory6Qhe0u9aRWqCy0tMEs1fz1JxIEK1DGvYWwj/rm6pT1GKa8LM1tERBAr3xZ1w+DC6TD66RQvn
KYhqRgln8rVo/3F4LvsMk32PBc7vU3mptaA5A057d6CNWu79yfgjCX4EhKV2p9gHvC5y33025/Om
MRnvWoYxIBA0BjQ9hKId3nC+GjmSs0yb7ty2AtHRAYqWQk7Mt1UEw8yz0oThwMsuffNcfXpNZqae
VqS2+vCJtVBuTV9lVKJRIQ2VUfZEYsjDRgjuh+WH/NFjivPRgeRJgWgz13LjcjAuF94zQg0ObvYI
acNaVnLsUfY/XK8qnZmrtMufMKocXS6icmzf1jv0uD8dEYSQU2qIVzkqMQrJ163TD0tO3HUskiii
LmXJEdx+QXcR3nTKtJPn9CxrDxJvAtiSzcWr1bDvS0IXwBtrP5w/qEsiEWzTDfCUZ60q0KCPSsep
ifirKRzZR9xGMjPcWV2zWwu5zDyANgd5gcFHv2xKBFxxI7j3YM3a7LnI9GF53GkTkMBHMApfZWwX
xq1/uurQ6rN+sO5W0X9junQ5bsEILkD1sC4u5Ax0Hb4eVRluRa9GLyaMs7SOqZN4tOV1iQda2c/J
baCuuZbvbz3+QAXF0YxCd2DtVwauAnz2S2R702h1xtGY+FRmU+g1qivuwO3WIpMoi2X7ZIpvBsKC
McupslYjj4pKsRTjR/rrfkg7VNqIgMYg2TuLNYNQ/HWPzp8esgIeAMUJhIf5561/iLt9cwGoGW1H
lm+GuWPg9xxLhrGK3RRE1tI7sQJj+Zhr3pFVE5nUT6r0Lov/qMHkIlDsJm71upAVsukt3DbVJG0/
lLW/o6UBN1PGcC5H+EGV3MnxF+EFpERqbTVefYQUamQsnGj638jLssbPzYBVt7gJyfLkQuFymeZS
gtCNhlUKFL0iaJ7RreeBEog6CQR4sFh+Xx0akxeEeKlMftFlkSWgxCRKi3FYBZNepcsoFwd1PJWC
ZWB0w8XDij/5/xLKAD3sAfW4iuEeFG1UTauI9yApWAAkcaxNwopEy9Ap0B4zF8JYQ8E/nMsR9j+6
2PAAncFa03FQAULZMPShfZiq2XR44z/YVDkoihpHlggoQ2r9IBi44vDnZGroxVOFCSAbkv6t934s
cPXvUk3WakYzrrlg5o5OKpWuqk/KwzpEjdLOHe2EFG4vomm+3AsMOj32lm4ynQzF1OYrFEtLDHKx
HX4tYwSnOA8TxVT2r7ISaH+Dn+Bm4bjjWQ/HYWZhdXpDkNqSsg0FhOvBfb310DtH9JEROJUr6YEr
xN8K4nFCIewS0z9zO31YbtGqZLps3gAITv0gCJQ2oF2kg1WIvz+9+2NGRl4XOwXP+41LittBKOP3
PB2bYV4GRLm01DPOnMFbYZ3+qFOeWnEATCwxp2WWXkj3HuwYsiDiSW8JInQpEjYBO/0LKAbL4Mpr
R0ikeEzSL2QnHQlBxPdHHwJzX47877u4Vb3YHHWvPdjaDWh2ypc1LQwhBnCHlB9AzR/yokledOYG
AqStXjHxqYiRNQXn9fDU2CJPQMFUIx/nViwk3TFukjtGbSMWEVp+A19nsiUVlcIHpvgCxTEYlobS
b6fZBtXwO4xJ+KNQrpY7gj9cy1aT+owhVrluWT+NyV+3PzIZPrWR3fOaSoyC1Hag4uC/dp0O9e87
dctz2TkNFsy3YL0ebLc/D2c/0kwJitFBQkw3q0LI8h2OKm4vSOVcOraRW2PB56AeK8ds7ShrpeY5
3Dx5h4arerfoFJssZunOAOwiuZ14udbuBoYcaQ3wCgieQnhGAHy9F2zO+m2+qht2ajoJ+F5hCJxt
w/SypsjNzsH4rNjaPKVgNbCt5XTOVsZCKniSKj42q7R0LuVObI8i6TK0BidUqh2TLVQ1LqHsbhS7
AgsyX9+4DVMeUXk8G1oRtOjhn7VDsrV8MmU3gcZNdHuaJFZaB4sXXAzCJd/u5wLTA1vM2zys2Nn0
YT4cOD2CAd6rTK9H5zbu5bT5udMxgfv4HT/biiIjQTdIgGFkfBnaDgdvyYrUk79vWppAGItDtwnS
5d0fryd0lrufKoMoolwraLMsyzPaEop1q9rsFtdlea5l8qD4uPL11639eRFWpoR2C3vKB/Xx0lpr
px3ZNCtGWXKGI+oztRz0ZTkfX3c29T74sTzDTpxmyiWkE2T5s8rkzTcIJrllMf8rpd6tZfzj33Iy
P8N8bToPeKowZ5uKrNx8aXkLqXFxgvuMGJ3fqZzDyCT93+1bzA0MSq0WMzbb4H14j8yezY2oSPt1
vdLmSG9TSc3uNrDIM7QZV+fCPViBTOB7Wl6M86vk+V9qzAPmXnGDXDe0Qm9h9OVaq+ZqnQa8WNfo
7DiFbO+xnx4j8rQCS0ZmmFz7aJloTwZL8pEr46WmYkB5VThxdSWI6tuBVZTCyPGIVNXyQ/KBVmHy
ML+LDbBQxHjtNYuQAR5cUHN36KPqQ2QN1Bz7IhgrkUS5sSKYTs9O/rZS2/E7cl2BxDyKNwA8kNZO
ZYhx27gASkP9za0y9F7DYFDuj930V3+NHdumwbBQir46R6iXrUra9lxdAk4JKV33+G1dkOwJz5C0
5bv7dhHcTiIHU7bYHNNQNc+qoFVLbdImQ19nLACJv7T1dnBCVSeK2C55ZtJ8lekbgtwXjbEHIUvT
32ziMQnq7Oi8VSxTG+JFKp9G8DRbDdaAsBGbv1H8sKuyeA8QWT8rryLFk74kkAwnDGkpHPPE/jkW
lMfP5MTdJ3c1hOa5BZZlujzlF9ag8P6yOYdZKhCBY3okm6USevHroupZoW3HEenAxVhH/r5qOo35
7RiB0AbIjNbgj1axHWZm/adm6CYg3cuKlWJHmF/eRA38NiihjnE15c2Eo5b1y+g/dGDNtnDWzOPV
P68jiJxTyRqP7F/P7nTapOLxXGK8e/rJPwBCqdSklFasJFruQIqSYLwCpG4Suyl65xSFHaZnr50x
Crl9SRVP/VSN/0MY+efu2BNVLiRUNX5d31vxjLKLtYtJb6GUjSAjKlmaEhJbIk4UnLRRnGnUVIGv
IpE78jFwZFeJvgMcXEfMor5CVu+c4SOU7ucjiAZTPTGqqR1IRowMKhzk2rUlj5yWH+jLRotyGIil
Rsy7r7pKfJdG/kT+bS933mBqWGlU14AUG6mE8WeJ8dqSFQeW8a/tLfGKhS7N+91s8SBiUhmPlsNr
B5jgIsiiWP76j+2a61s/fqEqf3ZZY3O4IDuN54Yh8iTMmlDIGoPuHzh5QSFdHrhhXQCP3nAhzB5f
FmgqKziaPIUx1AhKzmLiJS9OSt2CWURMp8GTXEDmbXj/rYdtZkoe6Hs/6EP/Gh4SRdlYgbOYQnvx
NIuHS0/KKs5YuTiR5HV3UzbRTHr74xpFhl5cTIQ17SCMYau6UvR4hh86bMU8InFRCREXLRa8V5PC
sd4MoaUbfqsPwL2XsVpMujWN+2zofC1BgmKK/NjckiRuoSo88AIrM5hvRq4/V3CufLFcEu0LkC84
E7pN87Aaxxl3n1qjljZMS/ISfg67NKW+3x4/o1/mFUJhJ+1zt3peXsD3us4voSATEzGbibMSTKJk
0GEDRD9hznszICK5rC/p8avJCRTJMQyHte6fk5CkTvxSG9YGJeoVhz/Yddeyj4LnfVAsUZ3jd3fv
YrCjC1p1sf8qoOe4kNe4EwBf2eI4ZfeEUyJYACxh4a3Pmp3jVLdHzFDtViBU/82MHZDAsprlt0Md
Av+ijm7Aq64jSXt20/xFyFxFaDs6D81fGyrVpbay8AEtCDfaSmG+Mx6nC7Nc7QCLNnMcg1eiit36
C2aqo9do/TVlxUFY7cFPQ1BKRQ6SKCjAZ9IyBMghEFnf0GhuK57HHyYyrMn3nqN30wBpPWqHuvYR
Nt8aXv1LTTwD2ppcvLeeCUQY/LJPUOavbf2LQRBFEHN7rrZuKB4ohnCCRodOfr/xFhLwe4xdh83D
OnsOgZ9Tg6gSlps65MjZkeheqK1ZG93NOJEUzuIAOEs2TJM9yEeOURovPnAxRlETxeJDtVfGu3hc
TRuMIUYyJf7rkwK8kEEglCeSHXbN7QVl4d5d1/Tm1tV+zR1IxPmOQ0sCJYTR4RoW2DoRkf37YDqR
i3qA8le1RpmzEaIoBuaKDaldkJcrD1vgpWocDX8aKLueV/oJBqKVYpeKDW3nAPvLXE088Xlk2RRB
Vb5VadX6MoNSEth8gFqpAFDjz759ny2rG8GCFhRGMPZrlkiz4RMzGaNye3RYuNBatji++7muxPkt
A3t4QYsNJBivycd46Cgzn/pBJdW/xR3e4qNLwTCcHvqKhYPh6HBK0TnZP2Y2ySWklhEhiIhN4qku
c1jO+WM54CXfjNaB6xpzIwwZVnsWV5TbVK8fb/MjH7DScIiggiYhHRZVQ4qv2CnoUqbAeVJhG7nb
j7lic7/i8XPGqYoDekk/kbaRR9BlJUX/r1KLCaWBl4SfH2P9q8EsPM74U7PBF5qBJBkbZrgCX+Mt
SLk2nkp/B0/DjzKZAAZBChSaFvXw3SOmN5tTRjRhMgsqo21qfCXjEJBJDOPqZ7pMt4qh41NFqGyi
4fDWZldwOyx+CJ7KwFB7BBZHh5ODSVwaHzZGSMMGyvdLZlzjo1b+bGU+teVIdCg4lJo6RSsq5RSI
Fh9ARxe/wTpP2yyuvvyR6npda8rwvnSVjYf3gs7EpfeoqxB//xLIojkZ+Ru3T2IXtKZJ9RP4pedq
7FwhJXTX30lSdHceGYJJSIYMH4ZV2guonVB9wKCWaL5uL/hUWSB81xyFCkF4KKqsi4vkHO2eitBz
yPJyGvC5YVTLVrmYm4TxeUMFVZ6k6+ihxZmLAs9GogbfMHMB6PktcVUDCA3oA5KONwn/K2IQa5NW
WIPFtHao9o7OwEFuMKIjLXfN+DS56t9jP5OEg7NJUkAm5UXzIuvM3+PFcIhojZXN6qN1qem0j6lA
yke+pTz43wiW3lDA+lD7m4BBTbE82O5CMjgn1wPHvGEaSaNY5I2Y62EShOBCYSvz4kS7uAW4qTAU
Gh2BkmD2G7OQV6h9VTB8sFjfGpPH1ha5OltBMjfxhhx8emHSyDYUf36mTyVv61reQLHsNMZBzbgf
X0QfVM/ypcVpxubpVML5oTV9gSwLXkAqhr8ru/wKRbr1nk6Gr+8mWASNKgmBVXDw8VSnbt6N6rx5
eEWRiZM+inDimqdtvg09t1kpUKQ8SFgz82fJtvfFfMg/QidacDgFiqvLMO8Zg1VxQFtg9RHh7vj8
rstYiM2wIAg3zLy+05/81p+DduPdDyVQTz0gif/H31dt94X9KlW0fTEEcd+sKWUf8DD8ec7PfZy0
JKVkPG0EUYG0/OhP3DhJ51BWXXr6Lueho8KmZPVbeSSeZ/tAFe3YoVyQ3eQ846pTQ6WXmpJEIkTE
iB0jkdPm/Pf1UnD26Sus8RjqGzlKyiomHr+OYANHvWc9aJhploQNkIi3PxHi+8wogg+2sCrkX4cH
nd/F6eFXEfWwqBnZI90kl+0eB30H/9/Ysj24RfHWERqR5WmikHcceQa7eOkZ8B1WleiLQwAFeig0
7nzl2oW0rlIk/RMbsjYC/L0Gh8Iy2i8DjswIxSU60xkoZo/mylCcdQ9kLmfcpwVbbMK9bViyeJbo
Akr5EJc9GU3ZGo+G2UtYfigqggNIXddLjGh03x+PolUM0UGTKgX1PWalvjWib5ko36NgcA5UOAnT
y84Bs7PR8qR0W9QxWfW/FklchX/NSuQvLelhfcdRE2RUdepV3G3YPK2DKYmyR+MX3ED6iT+5OsYn
f/QH/G8/fDDooydtiQHWGn7QITCC+XESyDzXIEzg7lUZW7aeFOkojSOjBqWujqHezkNutSkiY3gZ
EcKbEhELLHfLqsXmZb8fEOhk137JLBesUnT6yX7OouLPb/8loL5r7+aUE9kwH/h0RnCKF2I6qPZM
d16ClFjeKBabjm6y/m/pHNgqyc9HD8/8MwpdKmX/PT2EMoozPA7UCh9ieZXfinnLVG/jEesV7w96
xD6oqzUDw8Xl69jmP6+o6pFyEmRbIjgr9OXrssCd937Zdt+ee6O00cAUXsj+x66neKYfCZz/7xT7
+KwswwyFHukdpT7JwmIJ06bUv8kAAF1sO3GDdbA3ucKJBI3b2JlKFXR0UvYJ+SZS9BTaVT7itpFP
3tA7jhTbyfTs5Zeu/9GLfaV8vYqg59eTAyNvQb/mbAosko2fKkJ6AL5qgk+h2CC3a20qQzXhOCh/
sBELQWIgm0lgZns36c0kILZz1YsXaCB28VYaacI5g3SrPesDFzGI0IZXWbrg2u22bVr5xyTHnoWO
iMQz83tyWcIS68ovRPKVJ9y0qLpPyAw7l2h5urDSBHMExBJk9aSrfCN5xwhoWDEFoHe6Os7q+aOf
muc4xUmiF8vaJC/WWp1zX/NQK42/WRyIojCKyIoM53JMCg9T9aQ5jjtc28bCXR4eaeDqXndb5BGd
RE1D/eyg7k7p3ZKKIL4BPC9YfzI1mtjd2M4vad67yLD8HmG9yqZeG4tvajC8Q9LomOzLGakJIN9+
Sogqd8/JFfEbhUIAoXMm3hGnYEydigu5ADgr3M12IEB16AXyiIdsrz0GpBfjlcPVZlxvHzPYgKou
CQ++aoRoCCNDv4TfchZXS8sEEtOAsnOu6E9Nc++AhIFUfqeBhTCb2sKs9qS1qjPBTJWwvj/a8Kky
Oqx1Hn8nL8UEjqgxdolLlks73nmA/WvgZb8CqFkOSIeItnTT6knf1r1oqDHi47esUb4EiPrJTPXU
WcLsCSJu4xJDrlJvK2DkupA31Q/nYaZDouWwNeFLzyNYBcF6+v6jgrVX1RedHVrxj1Vi7xgppsjo
UgBCMXInmzqPZb0a0IpXtS7pChg4V8X7RlYyivCIsZHyDFfOkDRRNVOzg7aVUgrHrMj8jSTIuwJ+
kIOZxbRe9GWbE2EfTlZuQ+7YC6Qur472JPJ512h+BTME5/SxGMT16NvN9RAhX/jtvG9GWMhLYzyF
3Kz8w2PChYYpFxdN2pTuUQYncWLLD+FOuMN/6jYP+ICG46EJVArnrkmdNbwMF7YgPtkljD2qtTeD
m1t16jNhbfw2DsX0hV3eY1ZvUph18x3CAoTxTqdx1bpbofSP3semaP+4upbVypvn+bm1Kekw2CoZ
e7YZUerhL9Q5CW8rrAYDqRZsYnzS+6iBYtrUZsZ8w95A95rU0VCnUa4Jknjc9h4G29RTYnRVFyV2
IEu+XwsvH+tkEoc7ylBQR0WYnbqdSGREcHzdU7Mrcq28zGqk/RzPJQ10SZYcLN/zPywmjluuleOj
Xi2jvNtzkEWD3e1LorpZvsjX479DLkxLHsOS+HOgq/bk9WE3hbmQ6fZnjSJXoeebldWgKMTt1RiJ
/O1R1eqN7tMY3nB1OqooWWe3P0MUP9w/OAuL9XZfDEgjxbjWKq6zR+3kOVnLBcoY9pmx+d6fbNcM
DT/hXzkRiNpsxso0peYQKeI5Yxjum1AcfA+9nJkcHXCOluhMnW+asQodPjJxsJL2IYtEhsTK0RYC
4D7WBWqJFTFNxm+ZWDHXKTidIqQ5y/YzP/C55LLGkSJg51jmoj9/Vc3RYTed2DSXK4haOBb0aHpW
FJLYJL8wvClXASe8Rsgh60efY3IPDJLJ1Rgwt4AYHRdxzPubY0X7vElg+OJPZlUSOpdynyVAYdoq
iOILJIfojiX0GiJZ58u+oQzhjGAzTgJBdnSl6pbWe3U9Ivvnt/Ddk3nmSTULNmR+Bfcku/QMsjVc
v+WVWaqjxmftyoKuWc7KUKZ2KL9IJoM7g3DhR/XFSR1IUCFLr8o6hu51sqauvDHRG3J0aw39WqvV
BVOzjrNsbKI2U2Qn7qEZOVM0BwbuzKdWYyxpu/cF57Z1dXhgBSf8BLufL9dijsfCYcz7TtlINJd3
PD6pVqpmca0+oEQceDMzGLxrvUbCj6vKJBwfvKRoB2QPYsbfYSdGQks9q7HPcTI0BFI2TUA8HsJz
sKnNBCnQxKC3STYYa9AdozuNLjGCPJg69SZhbnz2eX1qXo6vKvR6AV7Yy6AsvrNsLfYfQHA/Mzyq
jkGp3vnofZq3SLqzt+o2osy8oY+8HVfmYBEt8pp1ilZPSxP4GzKYFxevlsi1lIwpWhZF1Iq6/TkN
xevsk/WUI8E6ZaNQTbF36Zkcszvej1bLg0ZxfPePpqv9RYcvP9IWH+LdQ3jDjVPpWugKdpyQd0t4
l5UutMC48YQzV29aMdHcsW4X3XtYFhA+qmqSK6pZprROej6seljmVNg3MPy0MCcae0E+FpkeOyaY
yddlCmELtcLwBfwilh792Wlw2hFt8IHcfVlGuew1ts/+u/ITHqurLmSveMtKEVUwhg6FJgHH8qpx
eoZlHoG3WJHbnEeshTF2+/LUO54/TKvACuBGlXgpVjd9DvRPixT16mfcgLWuBu9lhEvCYVS/JrNl
5OYkwBS5p9F1I6d4P2N27QLCeKyZ+3XK59InLhXpVBOQHTRm1LeI+a7ZaaWiyw/CLvyWKdfh3ryy
t4YGVQ8m+JJRKFKDWGjCoXM689mx1rl4HxdjBhe0jnJdYtKpa2Q1kWjhdTJnkV4hKYMmuDK47InQ
Xg3Q1E6DO2yWv9wyRm7ausMEnluvL4+3CUCkW9bp2Bmzvo0CkXC6mo5o3GBXI1tTMfNUsYN0TotO
8MdtrG/NYAulgfSLZRVZyyL71QgdEpAgM+QZLZf1OBt0yMo6qSmsDQYsHFBXJtQRLAsY06LekmL6
jvR2gIiBzT58KmK6TOr1TtevIXgczdN+j030UkWL1lpW6RFUIfYj0qDHvO9Ym36LV2kP+N0EVxcv
GkHBSY/tE4xhEorChVCqaoAQlzOA2V/Wodmxvc8WvFAk5Zr2q4e4i/wI5lWC3MkzjGvCYNuTbn7C
pQvRnsHbDv4q4WEGG5c3yQM8JAJGeut4zlbHWGgSZX0TSxUZG5BzNMjVoZMllwsQa2lKTYeXVlyI
nshdaQ3oeqFb6PepXESp4B6GwPhgl5xq7m/y4dh3LCzlepClWafKoFryX61xXddl3HD5AMINEa7s
45D13vfpwEe2KGBvuGwxpVqTJxXNbgvkBoA5o/tMXHVAWtnFP/dkkc1cxc1m6S1IY2z8oP5HPWlC
WQC0KPL4UhKLGW375EYD/EsB3ejKJwU9pyZ71EhXYju3Ozm8BW4Kn/7xpQdaADZZT91GDmysUJDg
xm5BH0X7cUCNlm9WBhYkGEdCeR9W4M2pDQ/5PhTjdzcUfDd2RvR6En77lhICYWSraNuAZ2JalGOe
wJMDcOHfI9I9yAwH8AgKw7mC/tPq978MbwG8Ufy1Ecz6cNFFd+6sXV4X6U6tFgB/dbfE4mh4BAvg
zrCu8oqM6Q+9wwOyg7uLXVae2GmyKQXwCAmIqQg7UwMzv1m0CSRcpOG51EmiELQNzrw2s68qAaaf
7mFXJAWt3N4qpQW549su9Gsz/dU8SGj/ju04KLaumhafaz6FUtZXWr4T4peDke0+cvDewDhLHlH6
lfzfCx8EqMsSISDK9hZoIJqKzXW4U9AKo7TI+KbGo9kKpkfR1l23Oao/K+UyvhM0aBq4bNa19Dis
RbQ+vu4119vc2SDfnTvw46j6uVP5TMmp0gqodA71bNlAeB+/zyUbSN6TojRnh1bq6swgRlSy0+45
QWUIa1ZpWwf2maXmEZKqtPUnZPDDgdjfrkQkm2XsbjsZo9du0yf3Il2whqvZjDSTaLNJm6h1pyDv
so54l5IM5x75lzuHPB/qd6tj30xYS4OaP77m2/4WSsbfgw8zflSLhESQotcPgizmGtOMILNUJxvl
thlYS/zN1AdGBqGtlsU2FN3zcenAdrSYenifgzmPfGRuvTa+Neb0KWDlkwLw9IxQXQrIYVMhCJQ5
9rKPbGkRmxO+G5yiSfxEA/vHp1fIxKawkcL1EUhSotEnNEV04n6OB/LGySj2dzocc8RqA0cQp4lv
/q4bK4cJgFlr6gwFOT1BEDS5TFJNLIaa35qcSIkFy0abb7bsOYZ+IP61/0/4TGx2RX9ByLiT/Qw7
bJVrEE0Rw7zd9B5L1hIKKvUjHHhXkcyCBpe8NoXOpOLIpHWLePKApXLnubfvVy/1HTY3B2BIfvZt
QlNpLz1mtQlF+o1dHDeRqYl3Np7bdOrI/aozjNyI50pdFKSdNDcXgh2TJnCAMas70Jn6hrxlVgeA
+Bv8MyhB/BdgGdVD5YWIrH/5nBqeSBK3ZhxfvyJDyFuebrALNj/KobuaJC/ZrX2uj/Fm553Enqu9
YRSFAUL6QKD/eOF/EehrrIe11Si8HX34hP6Bx3ZvJAKZZDl43S+P1hENT78xw5hM82gcfkjDQCs2
W76UWgJolmh9uONPMx6O0AIrvUuVofc93qArWHtS+qlbjrfyD5XF4rr6b1NSLIGDTM5c43ZJYYYe
CegQUU2lvIZ8uwt9Lcl0Mo/kaM90U6GlgdDYrBtIuIz+eQqpy9rc6QzoOcIDyRDyU7Ex1CcXRnEF
XGGM1fePAGLZ8BPOBQd8VNWyJjRUjTd6PjEky1aAAxtgTR+/bnKmfaU883IlTE8Ci1NgWTEy4ZUZ
/SgAM4Gf6xxcVivgFErURQV6BNXsTH56zG3wh2br3RHe7dmoRxM1GSLj56zi9KNSuP1OaS0GJNWQ
ym6vZzKZfCDEfkdIUma01CUjg+Geuj0367qMV9lQmtakK4IE8Ze6HY1/tV5xNeDjmfaa/XMCER/Z
8YKUHp2LYVPsYpVDg4G4lzWMuUIu9K/NLP3dTOKA+hk9azqPpRNciG1e7vn3Z2DtwmZkrspaAoWX
lcS6XN557AzS6LSnrIyy3qu63C7q8QwATX11Fp+kSOYO2s3HFor4mfu3YstPmdTDfUuGhMbF5Bq2
1bNhh7y+u7TZhDLmtZPt3R12Me7PACXKtpV/C8ZZZU8TvSBIEkUBsv08kzWuOs4z/dpRJ7l5Zary
MJ3wl4XKPV0hFk735vi19WjpeRfE0Pzza5lW/o5p5XoDCOrJ4HdkoA2hMXH83czgS6DRyuHH+rhk
srXDU1eSeRMj6t58xmMZYQeJmhEgqA4vPMI5Nl5WSlOnUIwHZeTKE1d9gE6mV+I7M5es7FllhOMy
zgjoE0KvQyLn8sLGfqYPfPVFqtqHAWbWD+PpSKVVhBGDjFk9eZN+/xWqIVHBbh5uCgIrCTSbX7Pt
iJ012EWx1tPxnXKbShQ+TsmN+Osw/4StGaLzp0MHvCLylxfGyjh/q8LJp4IYa15NI8NrGBMQeU/C
ujcvltdoynCi0K39M23tBqvochJElLUGjHvAsSwIRJeoUMZYvgVthljmEc4tEbWeGOFVwNUMxGms
o+8eFbD3Z3FyNSDPzzcI9AuCyeVgF8XH28EM5bk5kPWYtQBD3jfTrELzTaLiyoJ93mh5+mJFdj6H
nfbDsjVuygdsv8QsVL4uVqLIVwoem8LnmWIKcDY0BWjWJLD6t45QclAIVJ4agZDNQZM2ItHm/paV
ZD9LLpHxZjd4Exstv9Sie1PfMKvR3aAOIoehFJh6ZbMW7T8VQzORESzfwBtDGEKHdSPhFnsWdcFe
xCcivzQ99O3zssKATjYi6j/+2HBihpQy1WKpbFiMpoj0Y1dZmp29xrpSCzC0YG2mjCZSSOWRc39X
KRCoRZrGsIOkPAWQLxZkmuJuumuIA3Vlc4Iw7F9CViFC4dBeZlJ+Z3iqbWSRJTdmnGMrqBb3LkG+
n4ZHHu64fTms+iJK0uov1wCYLGWaoHoCKjayDDnnO5uwEXKXoApbUP9hR6Oe355FWwvwdmd0D3l/
dgYnxGQunghakSp6sSKp1ryYLuJKwTbRzZGJ9RgLW3dDzBGg4N6FStu4im6RRHE9SLz71ChrvPav
2YzBIhi6g17lJ53Cw2/53bKj/GyY7Lm9Z35pddRBMaIIpPGi6zrL68k7bkjK58QWuYj+idgLDRwf
8nATNxPbnSahl4ZRUE+12Aqsxobg7H/TFabK3ZY/FpgzNW4IdJ8BXMphsI3vpR6UwtfFg2+xNJ/T
2L53Hsw5ItC5BdR+AH7xDlZpLuSTWU0zyZtCi8lWoVQVd10qIDxGtLPgkFt77Cz9VA1EKnUcQ/dk
UhOSTlZfmH3fI3ygmUzzc2Y97dBMcr2Nub/v9rP7Ko7F8SOORby6aIfdWi6WIuVfXE19blVyjrA4
13zy/0+c0vRwmeRUMiZhr4G1Q2exPHSNlBBLyEWEnspO5GGb393H5HTsxrjkqmXHa+kqYtF7vpqS
ZLXF1zMzCB0NkyRbHYUmFckzT6d4MYGWawkLEX2mP793QGP1TaUFiWkTb1jXv+kuhPLZM3h5ZM05
ukoiL8moRiAL13XNaXynmCurgJkAw1glHzr0dWlEvtQ1msX2Ci4SWcsXvQgr9iLN6Gkxofxl/AeI
gOLBFnVI/I1KL+7ialowPSGRAYpzhxns3Cy1vFl0IbOC9TcWTAeUXb5Izv2xDR4bJiLCLNRc2Izz
uOulM2ZN/v60ueRGwdPgAsfv+5lCOrZOYTMRFUJeBFqI0kL3Z5KQIxu8sT+9g8J5A4LzcyDglkJo
sLSUx0yBtnyLTuFpwoPZU2W5R1fEl6oWzHgZN6hi4QQ0OgZG/gf3pxQRyPWsU1ren0HfOXNQ3VRI
3KcHAnBK/fRVeLuODhFZ+rhUisB8noB36QaBikiS+jzQEztHpEDe39agpH+3N+lz0EvxgBHKsjnF
yx/S45vvM/r/E7dBvAJwWMG+RqnIAgPyS7O9Je1Q+neQvwn2Uz+9c2kbBk2WkghUppvRv/DXFLHt
gz8q7J7CXIHQbkGo40/nGE5IolP0gqv+y2NFOzC27+D115YwPz53yYyd5HmumqX9OsnVyugbly2R
aJUTpYy6D8SavND6CIBPuBph9tMPHHYDGx0gwO4J7+/XRZctWfg5VMCAE8GmkKZCTYm/0fWSTIQm
8WuYN0ukQQGNqMJ7t9dq/nB+OCnfvNAQo6/pbF0iD9KAncCYonA+ShxCgZ4+gmBwuHx8NcHQRz96
XYEkF0xeDG2NmiuIc50GNizNAGqcO9mgrDd4DBTlUnbR8D3Nej06LPAO0+RhOZbIau3wiEBdrLVc
eWJeICEDvZ+4y/qOjajbVbaV38Cqj/hwX7vi55ieSlyEfwOxfWpYEv2HKsfjPZEiCZd9P8R/7pOH
jqYug2H1LQi++ayIdw3XwHbiEWCOZ6iLBuyuolFJMwDIov2RMdkLN9Bc6+g709O3kjPkSxbGGRZq
GV0LhetPnydN7vHprlg6LLnO4/V/f8zGO30Qj+20QQe7fCVcJ3z1kTsUMGkKUqyn53JTM7pp4Vbk
BxlH2oeUfTJBgQnViYiEhslH40mgQoJ2iqPqwFEzk7oqPOHXnGTbdQEvbir5uuA52V5hv/1jH14d
WSdjM1BYy2/UpMr38CoYERpfS/eXve0mp8/UP7C3mPR50+dQCF5LzKJeT+XHmG8uknWUWjtoUi0b
qEV89nSTuFncp9ZzRPgk+QZ6S8byBsA0IcEk/hKORk46BE/ClOiPOjBO9Z6MVqJEeyksC7uPw44Z
FJDeB+4KI+Jdq2WY86rv3AwfDSncydyeohDDIHNDXwHSdGw50/NA8JZe/pa/OgWchDRcjx1x/wyj
wXJbYNzg7U2LmAAdvblqbqGZPQZ0HBgtvMu/x/uyChOvciTAiMuPprn37rOw/xRZhpYGsZWjiFrt
TIUJSXHVB4Fw3tgd2ktQspbEJF1EDXrnFz1Kf2ymPCBIIpNrMl0M+znESK1S+oJPqCovA37OKqI7
a6rSMU1gJ0O4S7VFGdObgczwhHywyQO4Y9u7gkoCx1KCEsfEHA03ZdVcazJX9c+M2D0qCYmlCzHJ
qo0Ae4l7uX9RNtFJgZs5767ZNM++NVGDLrESuwtFR1mT2U3cR91IW3qukEBHXJIDbk+s5ks1eu+/
BWqB6psRLPbE4ug6pDaKR38Q+Bkhkt7m98M4kMekNSLFfVuXRfFz3ccs5ltEms7yfXJc7TKjW3Ih
U3rB1UTuFbNh8OxIYWuvBvqpgsiBFGAwzZchAns278MrM0gBPRI2jxnrrIRop7/zIAVF1RQS+5Dz
jOxfJsL34w/ZSFxjBxMPtTn9lRuRw44hQjuIStLb/aae5X+4r2OoIzCot+nBk1+v+HFJvenHwDqr
Z5/jQIoSbir+p+h4xXQVE07UBo73PeEYzudhh5Z4Dv1AmxFepN5ndKfbYZIN6Y/9HYvas3+zbv6s
U+6GK7JTlqb4SS1g1ZWNHVx4VWp0A1Eil8RTwhm8tB811ZvXNiw6CuJNRDtILkW676dh1WujaLnM
Mt9hnlkMHtXhWo4uZo8nH41QJ+NjPyYZqHjz54Rqce+XO0EnR7FmIzbpdkj+3dyytIuJFqNcbc/G
dtlBf/piDbfXJJIJ7hbk0IVFgSC2pXsWPUx76LIRcvueH+DV7UPOoYylaB8cfP3AQBnUD3PNahjf
vqqAZpB9AXVQrOmeME8/JBy4GO5C5qAeYLJCya8aVAAvx31cRScRifWW+9iyA7Pm+1Ii5U1ucCrq
1IShw6fIUhRGGzIOArAXIdtHjaVrI9psjndNZeD0jDW8HDjuSLznpcAJ2VZ06Htxk2EfvpoNfINU
RcIZXaS35mqLXd1WvuwCBijWfHQfeSiidbS3PsOvk3UQFllRWal4KBgLTqDq0fY4wJ2G1SjbqNej
WqCDAwxBpcGQ2StIgqDhe7pgjcqPI/o3tY9Z7ks4SBwBmHtltjNa/usoSx5LAUhDZM6TFC1LfD4F
fdpbVhd6saa+YVWAD2Vs8nT1mWG6hBVrv8RMgZ3vS+YyXp/6SITUlxSVuXxHjfEhWYwleL7T9PcE
UArCrb2FkptGm9qQiLrOXIV+JlOuEkrANocp2NhY6dzfheJmnwGSk253cvD6jpeBHCM5yAQWYDz+
WyrFnnecxKgrb5o2aqvf+hh5gA1u+WbOYC3N/AoLOTsFNUasGQUxjzpvn6wMi9tHPZkAssIJ63Q1
yN3u3cS3uInKe/ARuz2caDpw/26sEVwqfnK1xgP4cSH+U8sv5yswH5lce2vnZh/aZjZRGNPNqc90
tMR5erw4GOgqK/zp68OciSH5OkHablZ2YUunGN8V5J2NAvJskJzZPzSX41bkFN6gxi/1aEDF+GG5
SNslB721pHDJTnHLNHVISh3+/CspddkzItfcueqG3ccKLwx3pgx9UaAd6zfc7qg3jeKA5jLg9spA
qdapSFdGVfNvfSKbPw0nzmJDA7eJ1s1d3O/CN36QW0M9vTcOFU48h0GShnux3IZ1RddtcdqhB++7
drRFhz22ZF3aL3uVDSzyDwLJpFpQrieZk5Cf6YE5ZXtMiF6O5WrHvt9ZcMGDrOkkYZU8BF+XEkUR
qrj0JOYMXqCSUyBmiqa3mq2sNIFRLXmPbStO5KmlsQNbZ9tfqHKQCyZ0RLXkgRR7i5bGZ0ZBh1pM
ahjZoZDxzzrtse6T/XMtjzSmgpIV5GdyspUTBer60cmar8RzF9qM84zPT7WU/9SJkRDzVq/Pmuu2
rK+BjARsphV/Mkcpiw+3LehzRZcH9p0mlxaFYhCBiJyCnE87dK/QjLstOHGiD324q+3IjAy1lrd4
sI2AzTxKysjqyESUyGthymJVSD+tQEX7UHqRFf70MMj8ji3Y2dlahh/5n4Xw/XWx7uE9wooUMuDX
LHAaIL2ynocpLoNux+N/NP+o8uPunQf+R0PuXyXuBeKNCon7QgSPY7ZwVOo+zK1ZfmzXSjjRxr+z
3ixmbJi2AFcF3b424g4JwveWRoL1OymULgIncumYf9Ct5eiL1OwqKqBs+VJklWL8L3fRN38H5H+j
DhbD0RRsD134MHwt+dcFNkwZv7Udqx+SjfDIRiEzCtnF/M1XXyrx3YOb3kmg4/52Z5c7itNu18hS
QU/dyAQ81iuENFnoNGsAgIVasb6dyv3kXLvB6LrnDlaXAbsFgTYWKnmkJRN8DPC3WUiJ9p196+Js
KYiyIqNtnhWELSyq710QMF3XM7RupzrGdKY1917oq8Ia7Wnnt9ADLKsr0zPd+PHmH0ovZCbjBRr2
xwoKRKcj/DWibV/ScnJ5HVuQ/rU89Xtd208eXMNZ7R7AZPZ+PBKnXIOj28GzCg8SHCTJ96k7psIN
1zCxkTPHk/Pm4E2git/7ehXukRE2gYeIM+DZy6tw3g7tVI1o8phq3VA6a3n2hr8Lu4V5/+jraN8K
sVQJqUu2kbKUCxNr68KB9bvasBC4ptFf0rtiKjAsVYmHxiteyBqYtoPfoeaYlOgQivo73+6hOMOG
80MOaHLf+pOrg2ZWDkP1Yh4Smww067TPyHK5HgQoUbFfJzXOhTQU+vxQ8tPEef6Zc/Dt8BiH0vGq
lQn4KxilYof6m9n0oXO7OxNwrNuEQT6eRA+GGsaNhvh7/oNQQRjBfgw0wGbCMnrrg05ar2Xg0a11
+mzTi+s2r3yKvky0uxFv7DocHKt8UVJYMyPmmYWUXfQoyXJ/yvdCSxmdxqZfZJ3+0q3d6TO/ZuX2
HcQ2PiVgwM9hBkB5wmh2Nn5JXVZcNB9t1T4b160ifk7VP6SIkduR9p5QQHB22DzOdeoWh/RX00PI
ihMiLDd3NQvoflpuYjEfOSlfLbVeXTkFPeIVomMIQiarKYEiAV7MV/d9I7GUJ6RtpDz1Dt4wJSHn
jO3TyI0gbg+ZN6kOr8X1Z3sDas89A5EVjp7HoqDnx6xV2X9sMrAocTINbF0gdFNX/fYRzaotAyJD
8amrN+kmOqj2hgq6Ejz9siwuYfSC7U3l2qGO+8zSpYSriZiYH4R8tWjSRtQV6RrvFGd4yinBqzyC
DHZu+bgPSdLEdV3MpOaUZse6DWwklp9xAL0nAjUeoDqqRiCFXzwWimbxLJuradmKau9jmQYykJ2d
Tt0g1rR/DW8S3+gUS/aoQDMwypffKNUfhdzUo1Pls1sDvbu0VohInkS4UoJXDFD56xcPfZCuKI8u
ezRJ9oOUSPqvR0HZSTgoQRPP8WREPbbdIWRip0dCoCsmjeHu0fDOD42KKHpbsUjfJIMPj36sq2Du
Pr2bPHy3ttf6ihLzB45cjppE4Xpeqv8O9KA4eCl51nKoXcZOgFkPrlN3gBHQYSFBDCrithHcqk4N
LKku0nmnSxap3eSnx4Xth1S2r/QzpINWoN//lhgaUj+wCrQyDcqCsVpv3aoxGCxGCGUJUnLapQSM
Mhx5sFxcN4x5WbZr0dRKPKT4RDsRzibsX86ESUnE6qFj1O7ZIf1k097+i+EDmDBJUHi0AJ2y3Ujt
T5HTV7UAhAv8V8nXS4y0Ja9i+P/8aGo4aE4iCibl8FufiBGyT8MpIvVJWozuaRdNPOKQlUZf+4G9
GWuADBVuX1i13e7klCJrTGk57gCzJVNLp84XpIjVUi66m9bE6PuXvxZJQcQffXsIg74+fESa9+Sp
1b/bIGb1lqdlVIR7Bo5qnlSNiz/LQMk7hw2S8Z6VZQndBJ6ib7xoo/G7cS48fFZdmUo7hx9zynaD
oTr9TcbLCxGwD4LuYYGYvhpcAUm1lY7sHP49frONAgFatFK7NZKCpW4rvgS4bA/fVTq+9rqN7SLD
K0JcjnqoXM+hJjHv8q6m2dMJmVZaGcheegv9IioGoAudY2qh3ga5HuJ1+ZmOi35Otg8NFXCamT9d
xppofmeijkVMemNeD8hHAnogCrqVwzsmRH2smgXXydL7nxABoqZqJmDo/0n83g4b1CO6pqV4acro
dj+IWPf2PuBPSCU/aPeQXefBsO+K/wPTR2gOqQuVmfc6qCRnexJ3jwKbvZJMJ3hL/jo9Zyl5d70w
N/Fz1CfvDYlrblfEA+4bMLYj4NgtENbun03yvKf7DtdHwIEgk5eAQuAN0ApknUt0JTqThXRZojjC
K2cq2KwCWbt/MqOlheUYUJx1OrLn6ajGHpG7Iu7X20OhFIkS7CHfOiVN7kj4mpFqttotgM8c5Uzm
1SauhITOwCLQkQ5o+Sxf6VM7lj2oGgtPgkWEPcxslbJzpXTbdFsONs5GwZEhar53jSZHRQNZX/uX
Gwhk78ZtAYKd2Wjw30L1il9nzkLVe55wo7fXIcwWwfORsKydSCcqHuDWCOlmuFdU/qUUv6ZoCD1t
DkojGKgDz8A/FvfIEI05tX0essZ4F9UoyGJHNVFh8lEFJAp+Jng03jUjgUtAQovgckct0xxYTwt5
BV3iuzO9va8qpjNnj2ArBi+bF9fCOkjq1B149Nrl9ATioVqQb7zy26xRe8VrJMmumiQUM3JiSM1e
tN2mOpWy+NAppr4VONqyIoviIHSR369lwxzbeBAk6+mIeGEP4BvGYmO81qu3x6GxxlL3vyd77VhB
p0x80n30ght7HYXqnOwY24fIqFDCo+UpJXdFZfBFpQatmVasZjT++YUdbJ+UYhPQR1oXy6QA5BF/
ltBXndrGsBDnwSJF4GUn8+F7wMKmNDlmwCU4doYG4zkrDJL+dq8Ak497nI7DreJtGkkECTX5pfhJ
mp6km+hgRtKaw7tz8ROgo3RRTchIfHWTbCZaT4yIBBQ30BP64scyCLToYddUhJeSO481OJ//g95i
IjM3JJx/MXSTudrGmhYq80OYrVbRXEHZ2HM4WGIcZ6WWGb4ITR/bLc6hJqol8XN8TivZtlpRiDTz
9Nr/GzOP3nNRQQANZLlf1tLEmLReUFBm7eJH627vxgCMN5vCQ6QUAn5O3UfKh0GoDj73Yad0AnnC
CDQI0T+wJtRUNabNh125OaKmQOMDq7L0t650BtNCoU4PoX5bkfmvmiYsLZuvS3snLJ6q7bHotNTm
FT7GVO8bR3tzjtWJD/6+1V3fcn1xFAgvmbZIb3W6IqjrXpqh/B13tQz07TR2fHiF/q9xlpKlPTmC
GjjvHxSeteL73H24DfqgnPNqLH10ca8NXYdZ0j9IgLAPS5FMaceK6MQ1wNSJn4hcsAu/w3cROqPQ
0KpfnUAIt7pimG0Sq0N5G5jrkqvXTejN+kd23Io0FU7txhV2YQLTjwWBOTfKkEDBaTqN16Skk4RL
2Kf8k6mf8zDkepP/i67L0ZR3Ocq+M8yPspRkNglreaG6TC6+aSGWLZboRVvAZZscO86ZtFUNrV4m
h89+Pci9Kd4ErLz++652VAENFNSi/n7BzpFGNNl6J+7moYpvZwU8lc1mTCw1ANhsuor4E/DmDuWe
WSLElfWv9TaKKpTjP7aVXwvmyeQXyiaE8V2JCbzGh/IaaxUAVtI8X8gIPYQ39PCRt79sBDNpJTM7
jLKpjF3Pp5qVb9d7LJ0zy52NLG7SEiXLFJX+I4C9PmGgSgTtUaW8NouLz/1JznQeyHiDeN5FXN0S
IRC2lmaNdYg271C5yN1LkD3jccYm4t823twDxz7mTnipHyMXVE0UM8zA4Q2+JL5bE4lmvPzOyM4a
+TqJ6URNmHtPwvjUnvKN4tdRIeuY2CUl+wm0UgXr8RdovR+d7XJ9bu5232UDtHQZR94pwyBLBKrc
r7m5uCvqjFxCKCtC3imtus8z8J1SNAKz+hq+ylwBZJIgXOi/HzQGQUu5iDTbYxCLWLxoa9x7r2E3
ULNfRHtd7VthAfwGeiL9g4KGxtJX+u7HdAL7hEUIT6e2n16hj83Y4cNutSbkd3693VJlLiYMBCU0
RB2dPYNwM1i6xeW0mzFN6tTjRoK5V0vgejgNwl8HyTqrlVShULgJguqA9vseq7bY2L+YZZhiYkyb
JWn9miljE08nZ4GiuOij0njxjRz6revAiopEaUL5AY9Xnha76i6Yr4krgGnTxuzVayl8h5D1fLQs
Onx+wy1N8bxHoNPribz2r5v1C6EyHTGRt/h8H01XThtOjG86H79xjQLDQjbwGrMx0L7Ri1ir29S+
t/UEqe6Y/qnLRXiU7G4grYtLu+bfyUeMAKhcEQCvOLPWSvYHbs9lgYhTQyyi/8h7REX/N/JvsgVl
elmRgSeuM5qTUl7t/ebOM7zN7i+WlMNrn5EB8c7INqYJoi0+6QS3aYuktjtnguhjIz5a+psxkNhq
Ce+P28+T8n0w/dEq8892eIB7t2BFfCHLSI2J8YJGJ8+cSrzkMLRFAch3uycBokqeLxgNpefnr8pD
bvkjJVJk00yuA9CZ4C2j1wYodTfbE3n8r5i/xmmB+X4AQyVtd1rx1SlWMMptrXW42pOf7+EpXy0E
9tRJrkgJ0uRP9k6wImSqY79u2Qs40q3sj2g25fj2nJpY3PEXrgTCfT6pDyHc42ri3dFRk1ki0RTt
R4rqRE3n/LBtyxzBgjNCBYeHs25IBS/kcqjscek9UkMyaLoCTBjRcG/ZtXGSPmS+7Z89Y2S2LNML
9Te3pAm4XWLoq/sckCtdaatrErJsYVS93e8q7eqJoW+vCVdDwIhyEg+bw0CwfyyFn9qUBrnuf4VU
QYdDJIhM1V3SkZj6QFhe5TrXO7sjHE7Hnk9IYZvMlt+Ho1NoY9Ux0nFhtj6imitqgJXHcVxUtqKH
21qc1wz+PWFWQ8FdLMNxmA3cGYy2vcuvq95cdz4X+qhTFeLcUUfNDURA/r3bvXTJQuQVf5FDaeAD
9d65I8p+X6d8UY14gQJda296zFkjbq/5LXy4ERPhSFPt7DZg+Ot31C1nsvImYJBNbhg+uLrohKaO
8cOmLDdAtAi1g00SIP72iETneQDZreWXcUti7Qk/2jbKsj6cOT+GjS7p4qo2aC4jTvBRFAzJU9Jd
6ln+m8482S3gE7AapDbjv3CgWvpIxpvVSjxfHmmXWm1PgBpwjm4y+SkY43UuY5dqqdq9D4K0Nt8Z
nXI5yNOcWRJSBlg4mcmM90WNbvf7bSEep/fMYtX+wEWswSXjORFvw7v2fLBX0YubyR9wcECtJOp2
LlKGPoQkrWGP7TTYENbLCJ0l6gZ2UfzNFi6OXRBCNGx7upPGdPWHMyXBTNISuYpjRT+Ils/08rDj
uj3BugcP0HF5KWYjWOFYbwNAU2jvdtMSxyF2JqDPjH7Mnsg8ifa0LZkZFHvlHsT2BeERp0TmT3mV
wclySQV/L9q+U0C8+knD8nf0l2BfQs/wEGp6kyqOTgmoiteL5VjbC95iDXde1iHG6ywTPJmZUrax
WNbK7ObAtxnIEPihZOSyAIJ/Eb9NLILKZ46hW9JCiNkAbhBjed/snS9CaYqtIbcZFmSBcFQC3xLW
xFaIdCVm0f0lHtbSMmb9Fyh5wXU1jwpXvb2+CiEvq5Sofv1/VkOTX+Pu16YdMrEZ9eL1isVPEu8A
kW8isZPvSGvKOAl11z/AZh3XkTMO70aLFR0jwyU6gJIAk2QpAzBdlpVo4uM8Y8h0iNcKqn48JoSm
Ort9hdmwx5sDc3LLfvXUdABaKTHoeouBUGeaTUPaf9RUmvB5ALo1F7pHWf2XuGQ/oI2Hi0/ZlUdy
EmOSEXt+lpSwComlFgRgrS06DMJsYSpSIE41Vf+ZGQfT8CYmtb5BgOg9azJ6/7IEpon3T7frNuOE
0+1F1fWzp1UzYKsu/Hs9ZE+Y5/Kj7AFFOUZPq4pBeb6n++WXyTS+CZRvM5RcD+B/Yq0eS2kyXDZF
kPpFMFTpvr+S4YtIvgX9+9jREKFFbFpLdxwiW2436qjTv+dEJpm/+TZQnhx+DjDWhqXjG3PYx11L
2L7odKNQ3n4wBcgIBC/NGPhlKd7sYGFT9RybFVLEHFerp2M9EXYDXeoQkLtC6BspLkXaaS14rCG2
UfsBDI4gMkX6WsqO1OYeW5Gp7b+2v+FWsXfPrIHvdOcAACV46iHDkko3hNBRoNusrQDmynFS63dW
8Xxb1X18D9B2LvK/kcHP9TGY9o2tkfReFtvjdkjt1gN5GF6JQpCIdkrv2P5sdhggFRptxnqwbaYr
LFQMmKIeffDZ19x1sMkj18m/Ti/rkmaM/rIVXfnyTVh3CHLJtJPhLr8h2S8JHbbHIdKk0j96kXgv
yFiWy+89mT5xw4RYod/FAc+mSRWwKEdk2CEZbSvmtBVNfvY47yeEMgua1+EGhUEmUbyhCYVAjou2
32h76+Ictm7lFfBtetdjPUzZW6nruPIzod3gxlopMF7yT+EJNPJBFYbzrZdPw2+gYzBGJh4vmSBH
/kgFZEjYy/+85Xm18SfEbsPpGXEuas4L+9gCIBWhI1SmVmoUDEQFXszdN38N5GIkxm9W8gRpv2bD
RUf4XRROXGX1GLgUuSGGv9OkuAdZUTklJY5Tcd/l/mLxKtqTkyYHtyTaJlINk17mrzN0lZTEjUzb
20Ys8KNL6ytp0kZPBPcQUqp+zOo+nTRVFWqJIrIAoMr8HoY/+Shj4P8OFRw/eoFAkk4D1g4rZoDm
XRYzwqD1YWgaAUImCU0+KreW+SCTQBL6g/xgLMU5ThYqpk7eD/BUrsXWzwSYDtf6i1fnUPY9KdiT
ER3NyZAa/mPT9vXxKw/c0LvgXL1uj6WrX9vF/S46Vttlqwn3OZFFPu5d3I3sHWOrO+HmPZHrf+hu
ReuJC/S+hSP4ui2i8OjprRwDEETqL13DDviTnGFLrsb3UExIxbGglZ/pCAbqLOrNqb6Y8kDENvVn
80aOMheoSq7a2DbnvTu1B1nexgQxWv9nzymxqRTPeZqWdyAT4c0jXIdX7P+u+Q++kCwxaQhScA6H
pYgfWaShYsl+pAcdrGonl/ClIt/aEEsvZF40W0GLKW8IETnZMMP3Ov9uVqW5p8I+g0755EaQPOmB
q8UWNbYrIvskkUocvAZhgOo5h8G1Z//5Mk2Bn91CPXZnIeXVBNjGPPR0jS5Q3uKkYgmDN3A5Brzq
E+5D2Ck2cNyWA0PEWDyizph1PxpXWjbTRu7Xrh6yIEFrJuE07P80B0nRhRC6iVGMRlqOvbRSTun1
hlsRr7jKSWtf2PXm7OpkVga5XKqwvO8WKL9JvubPXoiuA7eYl35/DKWpg2EPcDguTCMcoeBbJ08Y
NYEuRLGMi1IHWK0mT8uq+0zHleQtCD8fTcapg2awdFIAI0IRu8WyX/twrywCDEG8Nimer5ej1dkw
MYBYPGblGbOF7OTwuKaUIUO9I1yQDYj9kE2S1B0N7YLQC4lLLTrMdCCYS2AxfT0c6jUo681DEfbL
seQSBpCgRV35nFXbv3v5hUcZ+FAGgqmXBgJUT0Sdf+3LZTKjaRWZ/pP8YCsXtiEsYFmlD/z8+BVO
1eiYZLMY0uFq/zHlK2IZmK57PR0LhK2QxXKdNbBN+eYn09YJEOK0A7hIRBZbH61hKpp8mgcL1Gyn
jAZa9AKAPKxiQi4UARWsOabRoroklvEpm/sJ6YuvKa5zQgPowDDgZDnPnWZs0C2O7TueWVTnorSp
pTBin1EBIsGY6xSZpRxbVQqQ26FFUIhK6g91KBfDdFx92EZ9JMO6k3lhGBXwCHJjTDw1MCaw1jxY
IwR4drTch1BhiOa/5dfq2wVU7LPMPxWx2nEyZ8LfewILNMQ5M1DhfcX+xRqDWvfvMU3BdRHYBP9u
cOOmJwGRm3duIc6e6OirTCgK1Qq+wKg8Q/OHdkZhTdf1S9r2dByVyUexlmNBaTivtMmdPsue5pM2
6q3iFlRh2pwpUC08tP3EaSz72w/k+VE+CJe9RWIcxvdhFtymQ650Ds0rQhpbjI5a47XLC9tX+QL9
FCIYn4yUg85MVxanV7NKhvzl77p9oUiB+g97gbAtt4/5uA9PrWC5c0YMsAbtF+4AIhdybVyNSpkb
us+Y3N18yi71bLSLa4eLgNh4jjGmN1MuVXzc3687F5DnL0tJtYQ46GsrH/V6OvIdSQ8pPyCYjmVl
HAnuFJ8CRKehlPiEZvCJ4oovAzbsC/DqGQytqIBq5KvYO+FDrpxmrOJJBH66PEOWHKkY0xaSN8hB
Jjk+eVIf6wI6IurOHxXced9BXB2ptshFvWxyclxhjyO6A9ikhGokFMpmwm/FgpaRI8gIRy3fwxC4
VrnfhO9Bpl98SrtWoQHSP0a1qc5yEw5jtoym7qU5GhqZ+6CpxMNGVdx+9npEQO9Dq8+u0/k4EBHa
/oaczbQwwAQXxZdPd9Bd6QeV5Vv/CqU8UbCU8kEnkzv6eBXVlQJg8TP275w0jwkRpF/bWGNhHLCA
KcNaHiehXqBXYXTaQGVxrT42iKCZ+DHOHMop34Ppaz0BaeV3HwkCl5xYCUdMkunD9ol+jhEwH0yQ
0tjoUgOajCB9pHLgDZL0FDYF+8SG4VE2OlNqM2cuLqttE1jKqPPp6yUjJXltYVd3wcu519QKLJR6
wgPXlkxB0RLi2L4ltOb6M3tXU9/Fr4s3+tc/Cjo/QZUcjjbigrfG9JsXT92y/ApsyUVeRXh4KxQb
t7q3bz/J1TNyQT+dWjPzEN/H+nd5Ddo/j1nJb5QPXwtPajZ3nPWKBOV3D6AXD67+xCumXj46Q2Jc
O+sCTjtMMHXziH8c/vEpXpcoKScx6yssCuYWGbiObCHAB0FUvAdyzROZNhn+ftnnz/eFYvHF/j2L
c2YyRLNJr1XsQfnRzfGsxQMx31FOdi8v2uHcmTS0rkCFLTdzWG7A35R8aBzfbDchE/mdzx6Pqyar
7aSvN/eJlTJWtoZsPiFMYLn6lZooJQ5SKhh/aJgbqq2DG76Oby13lSor2SEUw+gbXbGeNGlFZ8uc
D1ox0vLrOjtR/L+Le7cn5i7jnFc+vTrZ1lSLsOOnaOgvoFvdpQT0lVze0rBl/EhvGZKOG5LK3ARj
mQqnD+dtLS8IVk7jOjDQu1NYM+04E4GythU2+xXVQyQthFZ0ceOZU50bZLe6Eni4l9/meNXOiJGZ
WSYRxTExghbLgYQXAs/RNbmIU1AwCtK5bRp2+xSrXlNUzTy/advS5UtUwtvNKxWR8DKhTzys5gRY
DrKRfQTlXHHBOY/oO1Easc4lKcHr3ljNvzA739QRKuzvU07aHWzSOdzWiaKHP28kDkAnwNrahVXa
vx75TQyJnZCsS+KC7tgqVf3LGtZazTysyMNJpz7Kg5QW9/9995XEJduoYWCLirOTMle/HDR2k4Yd
ExQho/6tNe19CcBosaMIAyO0T6QgVWyItO9J7cX6pWqycr31k2xi5LXnpud6q97T4hHDllwpf4B+
E8vpMolubgwFkI0n2gk1WncNzC7RGfVOruzMd+7CGLNCkAAhIexqie95M1F2A/RSa9YHrq/ZbWko
I5iM+DiAjO97ZftdUPbh2ezFokKW4y30IG5LsDD13qajN8HTQ9uscdbaYVUMqNUseObyk+H/q9FX
/snS/z1rHSSB56Z2NFGiS1/U7laCfxA4NjNMGB8fJ+ZZisj9Z5FJUkzXYjqoV+DFPty/FoBKaRMq
yDxI0RnE0lFXbM4SfmC8lUL8BoB0Y3gxSLV4cycb8X+NPqlxWS6mDnnxwnofQEB2d5pXkJrgfYa7
at5XakR+LY3V4NZKCDpu2/i+8WWkm2sukpkgrf5dX65f9qLYgu7mE4LZ3PKWSlXpmv5IXHUQMIE/
10MKuwb91j86Y7mg5LBmdTTQmUqrbu5qmhN8E+d8d6jz3N+wFXbLZooD7n8LjLdPguyAPI8xayIO
cZyGF/nhnIGz6DppECZbYDX6Ct5CcasoGv8nNkpD1NPRm3KeaHaXSyMBEojQwky3qCydwRMcllUF
uLJvRUn5N7G6bw2ChMYIb08AW1WI5F+yoomLHhHjLRVugYhBec+FaUF60sLYv0pUtyaoN0kNFNWj
R70uRIVbYcYNNvRoYjwjxyBNhLihAZ5sIFNofuVW6hzfqhJ8zscl9ODOI2FKK3acBUW3BVfgljmZ
m6jrsx6fBmnMwrr7CzweuZ8E3FTZa0sEOd0vZLnUYWubAGEQgxipNPZlEJr+HJQKLsMArRrV///t
oPSCFCWbKvgRtYMIhGD7fVrPcUtvxsBq+qaKWZSgznS9tcXHunLQnocWgaU79YLFJ20/g/qmSn0y
XxSLAqOSCxiwYgNpzZpsj7xPNmOhsxF0zmuNG8iIjLLJqRjduTd3bVESwyl6X8Q+N72PmiZpmhhk
fUlB+nBNd8JJe/U/afYzqAtcrYePDf/V6x9KOpXBPuO5ejahU1PpamSLCdfUgFLWNAr7Puulu89I
hbCMqeNnEEKvAbfPzkSBcPILncCX39aFmguhN1gVIpMTtqUyMamqCQLYDiEwjW1okoHaiJvFCsMu
C7TZMiLKn6Ap442e4l0vUYKgm5SbqwS3Wfy7t7trTUygDt3dAiA/ogoT9VADKze6u5RkLU9Kidkk
vmEHhU9S06KRlYmOv6W1yDquQm0fu8+JaJ0mMwwTIcIgcfxdoeuMs/UII2B8PIoD89zH0ZnZgYEm
jVfFHlfVnPAcr4RdulvIv9gERCG98ynzqfjbmLi95dSdARBw/pVZlHQF7qOyVotp5VTr62/MAlkt
XrM2+6X4Kl/5Ytox5tHj56uF8NFCuosyDSVksP08nWwBav6mhrs9BT6WGhvz92V0c6kt+WsRuEVL
+9f95NOe4O3w6wml3zIKkAgs4Zi5MJZjKPfgYDzmrr+tkdEKsxt9c+xj2UXO3IzWeVdZzCWujeRH
GdTCI/MZJU6U6P3DMybm++OkQh0YduZeJlCgIw48lbRArO1q8WrBAIFPa5x5CkDYiAghF7SzFD9H
vBNbeO6ndq/DTzNZLS0ItarGk96R+/VcInZkzFoNdD7gf9M5AjmxHgBSFWSuQI/jD/jCNHuAaUiy
HX7kHoe44peFs8HQb50q6rPkKJmxrL2cCHNugRuuftzJJTAlGxVZnvBTIGf8tVE44nt8EO/bMNmx
9p92sP1hARoZUGrAlQDLaPXHlagpOzx69hjESfTjMuQlRK3SfDGDplQR5Mc+2hwwODv+uMvgxtTb
lOyTirSh6vFbbz7syf32bkWAI5uh0xQ1lgKiay6nCL/BkfZW3Afg7DE7Szc5H52JFqx7NnEaAy82
yKiTnaAabxqWBIuJiOj28bwWogGhVw19/X3sKXpybPfTHryOswZkesodh+MDaiczPaiNaizp7Mi6
6gLpCODyKDl5qxdmcR9IzmRRMmkQ2kiw4Exs97sFE68LHPx65AywnOYf7s///9gDp2o98LX6Bbsz
nZUURYhZ8ZNSVwikPIBy5HxLpm4gfYSU1SPIYRz9TlOc2VdkA2uUdrvQKXYSp5qFF+QS/iLKAo93
9MzDoumAq4kdh83DbMoH5LNFaIqRRTLIWX9OWwtKPN8LZTtgD5e+piLj3JeRiSh3dEMEGDZf58LS
tNe/3Ak7MWMHrNVYhJNho5cKyjnNBERYHKC2/eAOlLfmYfELKlcLW21hGgZjUvvaKnEEXZUNPN9I
EQVU7eMv+/dZ4Ln3ycALB1Mf0fod81e8XUxTx4Qn2r6+3QQ3P+KuELY3mtpKIP9oWQkipJD2PZDu
RNEus9fXCJVC5tAS5eZkHFjJaavYiqO0tOOCeLvD121+0BmtIJ2zNEOuTsHB2WFU349FtjRsVug1
p9GE8T3FYMalcZvQ1UxpIWodrwOF9BTOTUWH3PB7swQoW6c1x6Sqr8SeE26KzNNB96Skh5UZ55Jo
Kl2GFcqS94/ly1voFW4cbUrBrP+CSV8gpXwhyM1EoB5QIf7rXEOg02n+Z5D3l+3DwZqDdudVIM13
5orlUoiMYl6z8jxv/MAApMPuJoOW2PemHwe4Rtxzk5EB1NYX4+oYKWZgDYKn0NkyRVnpTxoYXoZi
B50fdcvj733hX9ejZr6fy8WKI8KKqNgIFczXnrkEDv+HcOaIdVRCRFlMWw7RAd5ddkHTWjVl220j
/qy+ZUc0/eTVeaHIaHwzFrHk6zZ32yRB2ZXai/ZUzDtB4PY+YPnZNJUiBwU8YvsthJ86RPhc83gM
iQo4RdKyY/apIuChvT9m1VAj+yTHNGtau5yybiCWh6hFREVVaYvBxvGtrlH1zAtYXUI+ItLUAYNS
Hxr7xow9Yy0tBZ2WgVfwwrIvbwKE6r+9OHftL55O1Jp9fSi26aCwo5vyP2FmwhMCnwVaXcSL0A7v
EUm3/qW3GssI3lYEwIlkqoyEWW08fjlA8Jb7rTKO8CKPYcD8XUAoIRBsUdqF/R/SphfkK4AiDntn
UZ4Xe/eCkvGVCxDCe1FWS1taH1GeS9D47D08gu9prGQkI/RwnjKnYYP2yHnLgLM7JO4h7yL+wLZ8
cV6ei0NyFAbSED1cy5fsjHMfmnZ6crkQ4LqU3qzKxMK0P4SnaQ8imyFEqmaHV3sAp1Z7F2d/6Sc3
It54uXZNNZ0Kt+JjVzzwQ0ehROgWotyNqhWRsm1o/Vra1TwzbMNGpTUxZe2RPys9nlihqdYSiKIV
ut5u8EWAzpWu3h8FxdPjsRBrUwsols45NUQZAiHh25cuJ1Bnr2MTHtuqKQwOtocISbbXfxV/lJyM
jLWHNIIE2ASudQzbFPfrTATxSCGfNtqrqqMY8+TRwGP48FbcoE/GAYhNqBLZp0CDydZLxJ2Dp9Q1
Nb3Tgt5Gyg9sQHMQ3VN6YJQeW7qaNqAyYF93jjCPdpjbGGszFh3PZCHVsJD88Ew0+GreJ7fWA7cn
lpWAqTWImDOIwYLjjQaKosKKl68tfZHvNAETkraGbWyL7rUta7efvFctJVv1OMAUohvHzKEWOe7X
En2Qk+9Wb0sys+VBw2zPGhJHIy4xJmHULLFCQOOg/2a/zGuB6i4oPx4b4F6M/ZCniRTNXZQ1uX7h
rTMv7ISkhPksupos96cZt9Hkf2jz8CjlUft3ExWQohaukFHxh2fn5dszx+DWKQAZZMJNsPEhOhcH
Y+yRdZCx70zkbguY4jbYPxSTay/TOgEUsRmgZQtmUxXwH4pyfiMWGoUBRGePEkgGLcuS9xUNVpyh
jRXFtDpDFdVx+Dd5/Xb/f2hRFlMfLJo9BkfWs+K4kYEyip1B3S9OfFDX1LF4HJda0M3R6zYBNN8w
CT28s/g9c6uIqzUp922IJmSFPjI9mBDoQs+4BI121DvEgX7NyU0PdiWmU/k8jMPfAWSfDJhuTxAt
AvSQG3q+ZAAD4cXe1cROewv1WINP+enMcpqnSV9vf005gJS8l+veBFFc/UYM25jEfU+eHw7IeROd
AYPSnqwzADSBWFQ45KOk9NA4vaJw9WsD8+oRQ+x8seZupO4ca4vZSsgrFOC5l7Cl+88TocvAKpiZ
11ALWBlb84TKVO8idm/orzNB3IKJiktSpbc4G8stf90pBh8QeN+/vdst4gpBB+P/Te8s+I+VlLkh
KLAfRoPv7h2bYCg3zjPyHw3VmOtU+8pCmTifdnbsBYpw3w/7vdp6AEhpvQh4CEhgv9koPU8jFr52
2G6tKWVHgQrBbItrw6rQI3uSvL+da1K7fJDIggmh/CWJ6AF0yuYdAd+rVhFWdteHccKD7qI9OYg3
UV2LPmQRDbLsw0001ycuxWVgU7+97wP6a+DnAn08KKvtdsiIEBp1Q5pY234puHZyHQL5n4qXpFaq
tJTXwMc7KyWrza3AhC3VG/GETTYc7u9eWLXauie/oA7MwBiQgA3+a9ycW3SFwQRUfp2X8FxeJpH0
w1MTB7RoVtOxB0p4At+thRse6TdTo35IMwOFj6WfbjdOZ1o0LlKBghKn3/MOsBFmKf8xfvGmu8XR
vaSxlW89uBZsRORuMce/GjOZlRo+wwLQSAwrgJg3+qUxuSKo0tjLeNJgaIkulezVwaP9VDrMbeJb
46xIpxaiHNuKdXVuwn1dGi+37N6rVR+oUkyCNmJouamemTEsDO5tGda0qPLjIixEQdZiKhUUEaEe
NCDLUqKb3oIbyS6TFQczp4jpjcz6fTB873cMggiGxn8pMAcNRpKJbdTlhGYrMnGOdiwyI03P4T6H
Scm454v/KbTpRzfyUbBAiqmkMgvK4omj3OGgWV6Og5uHIoqIcZL8Ga5o1/EVCtuf8fEKdVYx65Kd
MSH+YIAJJ4Y10rfw1zvdKsg2vGz9Yc8vrDm36CNl8Fz1eOxUy8SlwnxtKLXU2/94ED7Rk3rJs7A1
n0l0bpIhlrfifTsamxb6817zLtG1qtDI8zYRnqWf4eNW8CbhxrrWTmxtoOFDlR6MfN1dAJI7j6Yn
Au9rLv688tRMUpmUQl7PHPvhglJQax3XGuIY9p+q1qVh2TevXdz+jt1uCDq64z4Qz+hYfBKoJEGv
w+YVg2piMmAq4TO+PRAv31HeTE/Z135fWqafcq/xqKEnQ0N8Pssn85uHO5C0O1dANSTOGl/tvmud
A5T7oJRovyHpJFzQ1o7la8XwtmvcegWW0T+3YM2N578E9p7IMINCYqo4vZJ+17SqZMv3BH++6qZ5
RZqxOt7v6UNkAIgVBsKXgn7LHY9sVdtWldQwExWUsCDtnF0uEnxDnQ0fo3byZJhgh6UNlXv96J2L
02gH3WbWwRIcXoLdZ7Fi0rJiZEM/X2N0YqCWXOlwzX1lRkIKHXxw9PM49nMnj02Hj8sgGyqQ+85t
GLOjr7JzC/IazTYfjqEStOAsF+7tsPRWGXZZZ4rn0R+FyT6yhpzO2cb55llXgR0AJJtrhp3b5UGG
wKz4tB9Yx/qEFipi4cZ+ROoiZwyEiXvfek/Th/JKraLjmilqJ2HGaHN2R+O/CloPyhwgM8v6PCg2
P/VeKuQ4XCxOmSBzBmt2Izg156YqGDXf8vRvyPibDpjCwVDKWhrxdUtYoN7l+Zu3HmHXclWsLbnL
GdoVeGeIYyVarHGrZCYgkpIcLqqSvIweqatVsXUnQYIC1cPI7sk2vc+qO3n+Nkbj9DOWEe5IZWVC
uJAxKzrN5UOox8mD758BJ0CC6A8GsQ014E7lUIQJ2iPIMKj+yrvf7v6qOSeZIxhn6mfVLLTnri44
bpqpvtaZN4SVLsWtbbuirOGheIMqLkUDc/KvuBB+/zPtIkqzVxgziqEKGp6kzjjQc9xY0BAnR5X+
ZItTiUMyuByKYpYxu33r+js8gfHVMvq49TPdgi6Mu/3QMtQ6GCJMc4b2l7i7+3ysuJQ6lqsuWCz6
734QHDQ9zlaadfYw3Oo1+bQIMmGSmnEc/HbMhOrgkqUVTAZZtt8TqMLZ5iYm9Hv2oPGw99WHFaB8
f3yaQLDExP1cH9Pkk9iIr3I6c8eBRD8/RgFJX+TxhXd3tHGzypW3pC1Znfqx9W+3DCC2da5JEMHn
lgq6j+PKRe0Xb6Ys/13weTo/J/DFpjn4DG90rO7qmWXeI39MGRmOleedGUREu4FXij7TH7sAjTgG
1LKi8aVHfvPisDGgKVhYBHMonQAVuoMwDrc2QbXNvPvIGGPoNhb6k1l0SH9yalXEb/fRjkr4hNo2
s72AlYtPV2bgDYAu2dcTyrVvHPAU02rfJg8qgKaeDSJNHU6alCXw5LvKwblYzgO4x2ZwxnF3ntg6
XfG3MRm3GmJjPPh4rdyOyOHEZV8zDZzkEeCNZsfq9txNOJCloPDw5PRleJFQS5Qt6H4QBGv6VG0z
q51ydyl4fBpv/84Qyw8Ky2psOFp5S2tLiGwPNBgPrv3UvuRdFe86KiE8DANUqdR+NdnEhwuKT+aw
SRj4COaGRq+KV1cMwknPCaaBQ0HPXA93g0OqrHrc0mzMnyymEEu+l0tyOoO1mpGy50smNvXH3H4R
SqJRtqOqrQqglAwmsYvcTQCmWqXNLvmn9hp9qi6IDik/S/MCgwwsXQ+lirIoNPdxqgwwnGmdeDSy
JY7lXvtTsI/0AsCSa36c9zgyJizUupDrahlx5YhdMTmgRODq+RQS39Ob02+QiTx2X1UA1zOCKctn
CeWSfx7GNbeQxtvvTGwxEB89zlbtJDlGsnW1evjekxpVLaC7HyeYY94MkYsuoTEfoEcx0DxhDxat
hVGvY4uBrDozgEKE0IEAZLdIGD3jLWuhJmaGg1lKbwtqCOw+xZ2lem5vmLS2en7K+PVQwIGRh6j0
SgSIFfnz78LLfC/F3zDMi6qMXqC/3DLPRxAFKOgIRjoxdsjdpdI9CF5yE2CjwyV3llGJLDs+TIk8
P+xUA8Ghiy+ueBlBpJ2hQJjO7p1N0c5xUZrXONcyr7X5Y3kiyHHh7AtUgcKt2lnCRjSbAnptMXQV
idtjjDdL8SYZTkBukX2OqlLpCkxW553TSegrZpBG4QMB0lbkt1d1xqq8FDlaUkIQquXWfAEAGPq9
R7QKdMnZ79yE6oNjE0Teg16FyKQ3ILcIEm7HfAbjvbxXgh22AhedzmxPK8j/3TvMnc+zcrf1aZBs
d+TAZ9Z0tnKz1vInesCb4XRzeX4jKhpjxB3dBgYCMAGx98hZ/OBmzg+isVQcMGSG2gochOhf8Zep
ySp5kq2qj3JTLKGEVxZgGHDNcyBSGNX6Rwgn3ul5Bf36wOrqLRpaFLpky4X6UFOgz8jdKcH0vntg
Crd5GCT1tXg6DZdzFwtSjmbZWckGEfwrLto+95XXY0efHrO63o2Rw7ts2Sw9aEU7jqW3NqRfaF9a
hGOV8IqKkbFGyEfbUyqCLSVBCQziUPQoTapnKm9ff22dlsidQpKngZ9WfscLOXw2UeABDVRzEMKl
qOpK0cwXfEvVC4y65hbS7zKj4Z3vZju2vxpk3Os5v0xqPeFZbnZZ/C8gZE0Ok76x40jjf7WN+TZo
gwT56PgiK82UYUYYFbQahe/AWMUhauIhZbfPOs8Q2Y2WPvVnugo9Qh6nrClbNoJV6eSAPFpBKWvg
0yn+bF7q+b3sncmf5fCzt+z3YjiDcbuT9KVRI2OeEXuzeg75x0liFj0sP7ZRRh/RJkjpXPqo5MnF
s4fts4/RpbulOG2IerIwIMRC5lZyRefF0mlR3SBxGM7ENEFf6+lWQStSDP4SEv9QgO7B7pTC6g1J
Z2XYj+GGFGND+lE+sp4HskX0QCCesBEF/MTOKg8ouM7wHfz3dw9dZAMQryCMs6lNb7UyCs5Tk1Ls
dun3/Lk9xrk/yybHrfToald5EDgi29ZFJxsb6YeaQk1BipFyQylMk0x+rmPyp3ngwysq1ETbs6yX
ZzvhGlvsb8lpN3xqzXRJq6EgEsMY5Wot7dGqRLVJdcMgbz6NIilM8ma+xeSWUsAKwSKnVA/xatxW
mhmWWdLCj7740O6JINwqgAA+/4ol+8TD9yn3SzCLaGp+/rkgOZt3hucdmX/kDXQEwqaWpUCHgNFF
F42mO7oERih8hXReFFXrmujiLQoR1bBZO9EjtgBdimASdNX1kdyj9gGN5OarVj8enGZuBLLzCs1Y
IL6oTqUpvNUE16SCHCOjk0foPWPaeCtlrynzKQnDbMOY+dcw4XoTZ+m3df3AWEQDET1SrjR5Nev/
PjEglj8EvqEKykCa47BE3A9sVcSr1nnHEChykcAMmhUO/WlaYqhZYTEOIu0B9idrK3xLcK/GdLJD
kFUL4ZThf2iV9T8N6TeXmM1EtwqwxRVk1KXTxewE6ubdf1rMcx4MdtPN6/JJEfl578pDF/FhZ4wg
Ed1Mxfj+DYgA3a2ZG1T3P9Q69PqjTFU9FcwDYO9UMOtDagEZhWgDQ0l31AGpWjzqC1CeQ1GF1RoU
Bb+fIuIsEe1LKec9GghS14KbWa1v7QZIExQnMclNEUj93ozowPQXWdD7WYjdcITNYXsd55eu0xL4
O0Zc3pC2AJJ8OvW4Qcu4iFLvYWVqdA5wxaUbh6yp+mpBEDFahTqzj14nKOeGD891+DYaWbC4g7MV
QbUAnvJN0NylfYQvK5MWddnv4HdIBROdJfRf/2O3cjs2Ty6zRkhYH+lRW7EDzURGDPp3bMML8tN7
yfwBsJhET/H/Ck9x5ydosxxAyQgsQjSMIcXkirXsJN8KMj17GxpaA3s8NoEZT1a/GZi5LE1VFCv4
xa+XTTuhBNbau+g29dZDQJYFnxlkNgpP/QuwZvwQYItA12UbfHF2+ceG86HhfnKIHgGiOU7qudO3
1w+4Y9CZjuo9fs287njDwvw5aaYxpMpUfkw0HsjDqS97GUv9VC8bRo+aESkootjstRQSkpExjU1C
J4P7rboDZM5GQFrAtjnQtblodBAZdxt6ys1I4GfeEKsFHEeO8j3F00dCSBW7GEdu4R2/9wPPUyyr
y/mi0m7+nGD9A4w4vVGp2Fp2J0NSUDMwSMF3/LoEBJHg7Myroosv6bza5BFMdEwtYqv46iMF2/Hn
YcCrMlV0mrJKj8KcqjxNfrUiA+c/rkO6Iw013f7yjlYMzIH1Zw4BxlCcKI9vfaSFLO/6REBN6zES
DtkAgfccoYjQHhjRBQ2yDuSC7qDo1gWQpVIOVYb3Wip0N686L9YywRQDZWyIvgCeQfB6Tg9NkNgP
4bo5fklTZMVCRgbRdSPIKoHJn5xEnS3MXhK200K0FebAY5wSXfhMdsHb8Da8J77rgzaxcolqqUZT
KMzOC/sCR4IEIl07xotIJqYzCZcM/FPcV/c21qI8zywWsA8kiRbxIezccB5e2dsEgcPyrZN9w5dx
5Ej8rrwJ47diDHD08m4LifgfJKXM1UoKh64QRwtOF2UqOhmJ08KVvN0XXhGX8X/loUf+1D74fNhV
LH1uWqQDWbD4rehSQ8blbCL5Rv0earNO6XYLScVRe4Sk6iyfZ5PZum10x7GuULs/0JgLZAZVSlOx
YHgdrwk26fU5M5IAxOCR1K+bM4saOat+PrYY/8MTy272rgwq3cU1Sv7noIpOty3I1+q98gRU3VR7
J+sWcpymDjC0v07BY/E3tcqou5lnYIdCg+IfMtWIkGJBudn3X+nL2W1tPsokzAR3Nu8hYDTqbkDw
FrNet47w/XpswRJXr0FCZC5v53KfPKnezaPLmD+scGNESm8YxtEL1TUxc1XLx2iUMQm9HFOHENdL
x/eGkKrNnf+W2bt18G/BRx75DEMmUrNDugR1iRRJRVucrexb1O2F44QYviK2Z+19kudupMLTffFR
Zc/H3aTyI9EOtbp1Y5sW1J/O06CMlzOhc3h3Zi4RfwoU8Nmrh2GhLscPPzO+JEwj4HDy87TAgW9Y
0a8CjcjXspcMgbludQEIu8/wkin7sxhqJNeKvRhyulGq2cV9PNDlZ3UDcmHbTV0vZYVtdRCuaqBO
IsNku4Go/Ctkqh1gGTr0p7sOL+ef5iqP7El120lUAcMVSlXKrQ2zmdPi3nR48bGfaE+dtxP5r0vg
g0h7PRxZVq5WuH/pu9+2Q/RAf1F/Je7ix/lVNRwLq3+MvBFxJdpXTR3tarolqWif4wk1ci3cWSOG
KG6CPOszZrJ+kfbPwMx6CkMo/cP1ZmBZaAvnn949cdy/RwTOlabQbSSLvdXmk7M8MkaSnx6Gb+IS
JUhD/dVN4phGLWDffQ4Fnh6l3y0EqNqPXMrNH/lL3Av7vXBPqyb0G2FopBLl/GRdcaQNu3rq4CRW
wYZXImQpuZc85GnEVrllrlBt0GnYKeBgB59Mh7yy6cepYi17NdAacv6doEIIS7x5hmppLhvV3DbX
rvo0rlLR/+oLJGBX1jnHcBlAOOnpMHfzrO40vSZGkI1qnZ37EFgLjxgfCLGnCR8V3Ie04AMiQzBZ
dKhlWYHLEFj2VlyfVnHPAFUg9VFI4Cj5EOwhEFfbOHcpfv7kOn0Y+Up4o7N2WulSw1tPqGOZDl4C
vsM2mUVbdQKoPeiRtYc3Kxu5fQHyrc2k525mmsRfsXY7qO2gBl1Z7lmQcWwojAvCN5TnobeUAx2/
nfmbrbdCPCto3wn6nyGiN4WnbQ9o0Y6as2kY5+0OjtPDbpmf7cPfYb1FJ+QryHq5VAzy4XG0deAG
kjfPf0icsZ2rmB4YtAy7ZqPnw6xVdg1cmNTXE4bzwwBOmZTbqc6VsMxho6jJeTO7iAUTz58IDd47
8jfAVCjEZrvUFhq49R/GUPA4RKmcNIx8r0YEKEVPOvecxlzoxmXrE3DDb53djdZ1cW1xQ9RynhKU
kedV8noYohciEbPGK/Q8rDcJUCuwFVgJuMlnsKbvn3FHVfXnOyWiGqV3rSS+sNqcFN4AEJLj1JG9
ua9U0OfNjsdVjWVsxyUFs3aHSBEfb0x63HHt7WIc3J+V23FPyfY6OsPSlPLw93EhQjCjswaCLKvI
uIuy0nUC2QozI1uVNlORN2SjNnY+bhwiX6PVbmaD4aBy11/Ckz1vfsEjUDPI27iDmOPO+CaI6qXF
BmQiSwGzXni6axKGlCII+aCx5uEM7yNfcSyGSU0/I3pyBadvfopeM0jl8YFVOMpf+RhVRyHYqIrx
2CEcxXrzBmN72QaABrPL7nU0xq6eMEvJeJ0LXKKGQfK9CTPxy83A5sp8dGsOqCwAE3rTzp3RASPi
mJxRNePkoiCzp2TTPFs+a81YbPPVE50Jxk3eKOYShYuWjy/h34g1waExbPC2KG1R69jx2VJ6MhU6
2YByFvEGxyXCTx9qKpUjliEtwnsFFJKlP2WQc3ChOaQgNEqpfP5oUnTypI09m31i6vGetZwBus+Y
dZkevCYmVIQNbRaUJynL6SajdQmjyY6nvoBTuo2xu7YEcve+B+p3oNYZ9Q2t8d5DtDpM+7iHhOhW
C+zkX4Yu7f2uLx1PVCf1DG5B6JoC4PuAndEbzuB07w7meOyuOdCr50GLldbA6qprsh7DCfliyiny
jndNqpIXEz9M5ydD/lCxzEi2ovxvRwFgeQri+AJ+65N/boFwv/sDKt+9Zx+Wqfj/m/OKHVpteC33
wOKUGjYk5op9f+2YHukgHBYEOoJXD00UORdnGl97cmg+3CXNtp/AiyL+D2HfdyQ97YNCnuvINNuX
LKBGfUi4MG6OFb2q5B9KxD2K836c73qdtOiYfMbPBI1uF5Gz8PhgO8/wuZi8lrB/4uccafIC/hKw
kuzvvSTI1dAf4P0PdrFe1bIuikUKpMg2EQG7AKSmK+76ZsRRBo+i26QaZSOGfjRdba8d1AAI77mG
+K+0diyn6Pwk/62C+DJ+drIksQzQ4lqnNGnxTl0bIM3Re44iJovaBkjwo0xPKv3EIgSsgJ5vAoye
ZboPxSBAa5zr8TNOR62rwbD6/KPt+/9SuSAiBZaNzjdzwzyP3wiWQDUhR6jliBy41S+HlZXQJqVF
CW4yfIqedbfC2huvRTP5lvsRej/WHUTWiefBZc3MRRc2OiWqok/acXHo5o27Ciq5sb1S6+RiJLpm
hbFMhkIunzknubuZWZwQviImE1AvTT8blKKOqfCKvqu+wbZ5Kz4PVN4zylLqQ1Bz1+cfvinc45ZW
fQLDt58VIcptUGsybKg1hIdf0+1mx8hc83uCdGlfsVXVdgPaH6UEnE3Uj+GIF4tIOTVa79uyfeyd
Hq1GhCOhGi7Ib0HI7ypEmdyDUQxCVUjZJUy8Sfuc3qcsxLOECy8POkLZIUTSa+RkiqKKidlcyfBW
Y/PoCm1/sk8C+q7b2emdXCqWEkoSlBhguF+aRIfXJ5LPbosQbWfgktRyEas/jp/x8H+CBTno4V27
ZDAP7mQIHeKPnWwo/rTyBNVi6gSkVuW85n5xFnoDpEdLDgGjNvcnPe4OWXPmupZL/8bG/ohpl0tj
S0cDBdXD6F/y2MbSSVHE98VyKa+L/zw2Jh0a7PdT5RNE2F0QzV7uqIQsfeosrcGpRhSPC+0Z385u
uXVX+qmrqOSsMTmAiAt+cKwp7AmdBofXRydJTySKjAMe/jCagDxf6jXdtnkPcBhtefHB86ZFDJTb
4anmicvMkUp4sRZT83HSXWbNW2zNcX4i+UJT2i7Jkx7Fa4pYQ5JCvPvftgoZVXuiGL3xtIr1yRNg
ekToXI6+buZQkm3Eb/ZhqK5QgKcVaiJkO+5+mtttG3Z5n7utAGwK4NVA5N2kXjYtQbnU7ZORgYvs
+G2IuBGtsuX4xigzutWuwC4EaOJfx6xqedojJ31tTFqvZllJhFdRCGiXktha/tsvZwH4B9Hu/Xuc
bMEtAPtxXy5YAcJeG/1bEpIuWJDV9Yc6MJXPRq9U8iW4RYSEVa87z4djptR/u+mv6uto9aibgvHv
m0vEjLMxPuNVSMkkmstqxcFbtaVYiYwsXDqsPwae648GDRHVlhLMgKPIUHOkag3uc8lRY3auLuWc
41tIImx4JUgDMVwd70VajNst5OdQRR09YQ8cR5mvEE9RJZGeOVEa/z6w7+aKgKMD+AVaSp9Fg38+
9I8J1xMytLNnRTwZHRNdETfJ9UW44sdc7/OPD2jb7cUUAE29vVSaQQhrZEDkGORWic8Bl2njK5aj
PbNLyApcfly8nYpdNNIDhO0ugHNsJFEq3+NwV/CDeRl5dMHXKYiNUb3AaqWv9JqyMVouK57Qi3xF
DQbVMXE4A4qzWL9NmDlYZBPR2kUoRYjVmPBtFqtAtBL3JHk4eLryWIG5Z5gIvw/hUbj9TkKHptLi
Uce01EOBSKa2qDvmF8IjaZE5fxnIEdbNAx5v+fKST4uENCFzZ1kMH6G2JKixW+ddADHIZ3Rvsxcp
1M69+G5g9KFkkiWcQsZ6iR9DALD89srWn9McVLaO8APLeULstJmw5mrA8YocEwkFBWJXwxZHlFa5
nPUqm7uuy5seaSPwRxXpyeN/c/seET2vporUibCPtNIUDKTdrTRvnS3SuFAsYRirddk3ezgfReqq
k18XZtTrkMC0t8quI4LjJM/U3zX4nVKIyjf034LGbO74uecF9gHraVLsWVEDi7/O0ufUrFaD5yc3
BjrS1XOhMsXgou6Eo418z6C4XxIM7lY1NF4fLUO482m7AJEKIJJSae1BuKVPxBd8W5UXHuQTJFN/
dDJgMRTIs18/r7Skj4lgjfTXmW3uJZ0rwPjKCp5jAtw2CKvvx3vD2R0BOmgfHU03t/st5Bwd4Koq
2r8WQ3hojP2OiYHwdrjsKYV6XULsXrvVOOYo9gsE80r0vhjYTuZmp22Eq7Fvai25s+Oill72ZO5/
OXzUlaH4TQtgYBRrzN7KF6Ldm2n8UfQwo0/nFwywcKk+YpDNavxUboyXAok0NTzH17EoUHSJ8xTj
4GhBj+lSPPqiMRX0eXqDl42QcvaTyvh2lZTqhZX2xU2xUsKBU6ZTm1+2FAjlxitpf2+lxxB/juzt
zvh/fOblLxHH3VT3ZrLtkoXNyyVa+AAjj3HaFX5hncMj9A+5kK/fkd/iLpvVZTBcp5OwhYmE4pL4
/8z8PoQkXl0EwVBbiSXJBrYY+mpYPDyvmDKCYUxlObSTWdcvX+k41rmV0AwGqgxzLcwu54T2J/dS
ndtHY2fGfbWajdvWmNvag+FJHsnEb0Rbu9MgRYeSA9ZU44XK0hYW9X4vrBKLhrKcJ6tBNt8p+oJq
S8gVy7o2Kc0xvvSSIL/sERFnKFQms6JoRP9gBJ71L0+efpuhVNF8w2fccQXKvNREIMKqgTv79DiD
5FI0hyoUjXE8teIk1mOiDRO/TXHAL1EuBaAFBtUafVpCxiA/49U4PFHSjG7P9g8Xzl5DXNv4JNnN
YUemDLVXZfD7sI2zf929VjTrULwG8JOFj6FCrnacnohLTW56mhEK73kV39kcrB9p+16kVGAro858
otrbzXt2X3UPlQX3I8KMianO/icjgiWLNHp0xF5NQkeE5PoyCHYOeVFe1SghiWsFxfNrbXZ5GZqP
wGsDZkz4SNVnLrKo+yKh4qoy4MvInJ/Y2Mk0p3myCA0j8yD8WWAX7KPH6QoKbQmpIrJbPK4BTqq+
CwcYOKLBi7VqhqiEAYHWiwajzveyceTJT1F5fhTGY7ODyvJE4QJVvZ4MupFKSt+PXWLwwIauPmSc
5fdHBxQxibt0pUrNptO7puLMHhkwANJEWcZ+WdydsrfgFgATQp+5mOs3YgvMvPGrXD7vr+xll8EC
p+JaWnIlUW/XvNY4+Yr/vrUs+1OYDezvwHLjPcCjFTucOa04ZreQF2F+liITgG7oMuJh2awKHLj1
64yqljjVU7z0daqgoIAYifEM5fxMCUyg/qpoBNsDAbK5Zz8QzBDCEG7r402UadAyPO2OE/XtDBGS
Nv1UB+92Nqofu+Jkhghk0CoCxEPXRAdAIW2kG6nDooA1sl4Vrgfox7X38Nbze0XPm5xD4R5ouKvy
kZUpWCF34lp20QYlZIdomrgxuHN7WWWbf5VubDA7yffhiZAQue6+UzBC4T0WhpMy0qQkNMvqIz5p
QDAsAlvtz8AcYwbmqGisL1rNPfRk9ndRePDAgoKCdJT+Ld9kwRKSA7DfGoW121piqTe4DZrEhEva
jxcgJkGXr9LGXNsVxdf+ohumNRRrZ7TOl19Z5DCrY16cBzMg9qkNNLt+XCAohEEcPMfc6sgPyHWq
5wCKnXcukJr5FlUaVHvRh57D8Kk5Jis4jYPUmFnTPAXuENbCS5dQ5lwk4ABMWFnd28vzpT3iYbTI
6jJZNnJAl4OOJpVwSmNmYnqyevCMSGLR+ICw6lVhg5AjxGCJxAxeUI41Mbt1AxujW2Vt9HauVNAf
2FSTVB9CG8sKpVoeljKwP3I3PgBcbUxQR7DkmqUIxy+EcLOFtswg+kryqC4u+csWuitXo9rKDmDo
ba3lJt1McsKlUS9lfUUkUr3l1rjUt0gJvaPaECBRUnKFL+y/kIRhJhqDXCfNyUB12HwqUOPTZ+9h
ssNtVw5Qi8brylPmuD+VsgHbRSx6QJdw9arBSOlTNbwSrMEYaOUQgrEIARRdtd2N+J/ko/pRREou
Vn0UxeHn2UWTfIdV/EIhFkXYQsXUvcsSygNEBLArT7oV7JWmmF0du00ZfcFcu6oDp9y7gGzBw/v6
CywV2DeejvB6A1EUu6itys8yQGn+T64ifOr3GBI3arxW/Qb+KXP1HKgFl/DnmIAesfPsgZMITKr+
RN2Op5jsEE9FR7Ox0WORi38AnDHc1MXM6hdgCxu6y+8rz6lYuOJ9wMHXBUMsKRDHBbkpbs1okYiD
f+wIYvtvKnGOusXA/aIzM7kuwsJWISqPo6ic1hs1Zz/a20rMz7Shx+Td858odJT/Bc4SZeqm4i8a
imINfPCN7XLVMBNQ7zTSDr51zi3FOU8CMdhsTJDPUp9yhhp19CLoi18xUMZFgm32Pk0ORunE6CIZ
pQZbOtC3XtmZr9bBC/fLDyi53KsAT9QYewotHV38pY+MBlF9sjW8gBN/AwBX7Qd08FDGXd+pYoP2
8J5I9TJiOBfnT12aJr5AXTioKtoQ0S9BONkCvmCoPrRdr+RcleXUTXymbYdeVlzMZxHprxrIUsnw
WZIElDflSBzzJTCEftcgRCzF2oSjUgERzlZuU7V49OIGZ7UeivmiZAh3kMlQBqeFzNaATdFuOlZo
tQo0e4dtin1gZYxQTI/x77m2+iiFfNBxvIMO2wM+6Lt7Awgt4NW1F8UVPsQ5/RpDgrLGoqeiUwS0
R45jVxEveL5oAQ2792nc4+bGjKd5QhtYwyFL4u7Wtm6+iQmb2U2rCfHZfgrF8gdkHD6/dUi7B29U
kAmiEM0IUgxSH5VcJABOCndB24LVHBL7ENomnLIkZWT6XxyWCs0zPBpWE92wPW3QlE/CXaz0rQKC
6x/3uXflYTHwVyPJnDagxy988jEZZ287FeAyZ60QZnR/bmnDzRSpqkYCr9yRdNXcexoKr9WfeX5T
GaEuU64Qgal7BGKB7zt4prNAJ/f5eTh7AyPOIRmC5iOTDY5heoTnALADl2L6PybOeTqLMWkjaDDJ
NELuhCP5IS3DLs3I4BF9kCfWb7r2r9TGEPCxQaSMqui/nijE84ye5Tp3tY5PLe9A3kyMx5Dd0/6h
8kRUNzb+5Pz2Yck25WKu9md4ZZMK9vOUES49K10TKdzZhmg5GhuAqW+A8v/N6/Bji+7CL8KS4b9s
wglqQbGjmAsmASOTibcET96w78/qZ6OLvfIOZkQzWxAci9QgRbJkJrIYMd9Fir5k4VfY3bp9k1Cw
FxEizv1WXqu602B24uOMI9lemFz6+v9eGD9ZqW4QGUoYC9/Wfc3JtzIPaEpwafE4QISeL4wH2q7u
OOB2089leoEJLTf8F/gndhmOwfTa0xA03iUfJOrJzoS+oLqEc3QUH16iFAXZVR3e+kXiBHcaSUlL
evupUiWk1L/6cr35jOWNUW6uyfoFtB9ngkkIFq+mS9xBTN+X3L83SWz/3fe0hvFyz102NRZwneCQ
rQ+8EOyz5t4EwhEiBTUAZ35MfxRPhYRZ1fqXBicYyzp2b4RBdn7GFW9Mg8g7ymiYN0o6U3FSQuCX
pEnHm+lxPmhpacpVe49yEPbs9A8HWADNKQgqIa5Zmnov1E2MmQ7FLz9pisr5naeTSA6mOi/nbRno
DdcO/yIecyFVP9LbqY0Z2ctHLtnrvMdpo9iaW/lajnQLHguO7zjD4fiFZlRYuuRPe4OWAJRBkD9N
mWnQOIxivC2P4eYwzAcjymekXCTyPTMI+huWjJpbDPHY3pjVKrfMfW1ekY/2sUQtuNY56gyTq5/+
3foEeWT0MQCLJz7UVgJ8KBEDrkCZKv9zKdJ8OINlK00LTv+Kimw2JCA6GLZ0MA35P5RLjokJE+N2
hSmuTm4YqOPNqjaJTXKdsruCgU/nUWG7UBtdlh5dTtFYZXhLojCIGzbY2L8N2KjY2TdH2hg25s2r
DHv9hcfORo4GIkngedVrA9esspJa+oKW6PHgnvHofL7DuFa3D5v9lxRRx4c0qWFfsy2M/geeeFBa
bGMhTdtyukblha74WM9VMOmTcFiRFwy81icDdmWh2i6IUtmsmbD7aRO1eC9tFqgophcRN3xXxTFN
x1U8KwLxYvHNs1LPwmzEs5c3Cqb9oxcCNNSjt/Jhza2MM+lFQJDvTPocqIOwKYnWzJ+YAPFbja10
XfT5aaEdKubz2EVBVe21Ru/fg1t0xasOH78VYnqHQdVKpvZcZ8utTkVqlR2FR0BXWAuMC950DiOe
qtBKpA19FNEcB/kIYDY6/ynsIpha8Qla4g5/IZOaWY12UeD9h6xOw/WiENRpQqcAD5sR7FRgMsa3
oQ3tWzdaWH6JUZPdK5FLHM5K1BZCCOMm6ZaUUSsrPZBac+1xxrZJwOxMBb+Nn2W5/IgscH/NrfQE
WWXgjYlIpDj6oSNTqkTnBBf5eZae0mh95f9zgXecklpOK/nBBuDP8fB6uoIzC212CpUo1m+V6g8R
a7kUH39Y+jzYZR4sR2gPo6DrxWO4e3EqYp/OFBpMw2uVuHOjZuKjR23jqLs3IZCHoCPjtf8uQv3t
g5J1kfL3BaajZh0Z50Xu+KySQ6N5DsFRx4QJeX8td3K+LsaTp6Wjuoev4uXVVxB1KLaYZKIOlL4A
W1pXiscy3fGl0FssiUPH/ue4aiu1/YUZ8zSz1pSwy+uDRsyB2u2rGUk/xcGUvpCrTz3k3vIbt+tT
w2AIKuPyoz8C/WFfrKMx1MsL2fQ5D4Jz8eMzZod7MXnHGEMGOemp9R32N1RxbCHP7vGgOegHkcQO
rUjIZMEuwDkAOAbmGpPS0u203C4O9MaWqgEg5D2CjCzskMZZH20m5jZxKRiPlh3Dwtaa0MrZ7UM6
yieyVIavTd+l6iEoWjJWOTUwZA1K2+TqqFoBGmQogKJbpXaW0pXAZnulPPdh/zWZVEHvzVJTdzwh
fDsXKyEW8uxVDSpzu1kQ1YbfbCjp67hYc8D4nsQOSilyfMC/vVqChKqA7dTMcU5kmZr2Z1Pjy+5S
Xjoa4TWpwzjFAiU6W2JoZhFaf/jgG5O/e7/2vPl55xSSyP+UzjHyuyGhze388XuhCnPUMEHvmR+g
r7QD7i8109h6ErRBcT+jFgjMuQbGYMHljmKiaRI5oxcX0zjngOlBirRGW+YS6L9dcpvsW8xAL+8P
HjjAZ0tG8rIm4cOhlSyq8Ss348q5LBwA1aHROJuoH4gAjL+JbqMBMbGjP/2UsGGINoKSJYGDljdR
dqhJ55teL0pZulQ+WMwWvGdpkvS6JTow4hdBURDMacES3i489VLIy3G2b5da4wJD4cGtSDR4nWwD
xt71bFxTqGfrMNZN39JT62xVi/OIhePH601Fn8lrgCUe4giDdEPDeXdduTPSB3fKklNNP9jvw2B3
UH+u0xDGeCKR/P/J/SQMZmljvXtMOI2g0kv90DQw3jGY67zjlubQTYYhGVNjTHcwk2IUV5wmCloP
zuOkcnyyKxVXvpVA3HQxXplEEHQpWK83N2td1mThBQk0gGL27pRnFMyzqhfKZX9OkrUmj81Lz9Vh
Y/6OozNtwMyfKB7z3W6wrv6NAI6LeUh8wsquVpw/b4MICmxCKs860fZqWtCRO+9ymRSaZRE4FmaE
PtgYiVwcycLSTf7th0FL5U/LOiAcBo3yyymQi1KEIj9Dp1rCSQk+YKUcz9CXI5E4uZPx+BV2fDtc
Y8IHYL9eFqo6MHmUWkSRcF3Q++rhLmzGpAtrN3X299s8U03NGvLNss6TjBL/i5ip/He0ZHKx2urN
HO9QZqKco+XwM0rfbZKnv8pQPOGO77V/2aFZPzpTUrVK9u0xEQ1KFYxhdhfM3W7OPvDazkjw5FrN
uzwY4GkE7EtiqG9aMWc5QIeM370EH5LQRkLjw9inVJkLPln4nEj0gZuhKA6YvAw5e55amSJB6Yyx
t7I0HepfaL0fNES+48pQt45Dz1e/ff3MlEPk2FqvJ4htzSqq4TJJXKBPRmqYkRjKqe9M80nLoPbG
bOo2NL2GaAQREVk7IEG8OVEpV8ZWhq407do6DR/R/AuJtVewSpKDJta9ZRUU4IdeLMZVuzRW4Iig
ogCLCLoAQDfohdXkG3M+nR2+VO9mpL3tv0Ax2Y6BP1wPMFJ0xR5Y7atYPnI3DRBm9RnOTPXS3MGz
ZVKlDS3kRcycTalit/9IZoY35PKJxA9TX3yxp+nOstr57ytcWFpFC5Vbl4pslF6W9wKLFugSP4rP
98+IXYPwgAAtIlRtU/WkYgbiKxWhqHThJn38+B1s7eKfg26ZUMNVjloIuQWXGR7+SfWZJpsZgqGs
27Jf8QTToMop6KeYkJDjz173P2LvVJnj1VCwqSgBJvSiXPS7vypA38MOkS9kdazYak1Ki7z2QtfQ
8/UdEhTPkBLYjUgOGZUu0rR3JHd3VRoRMbdwR9oC55O4aqhT2kP9kNaqlXHS9gA/puNbU+A8PNei
63mQeeMoDzoSxxpHNJWX9zOZyHn0aPY6JICukytdFYCubtWhPWAAKkVwRIw8fc1i54p+OSWIYgWh
EIfDxJxRM1m+B1uudgzr6/ZTfAN4CtlXYbMRJMKOi3PJAmrkZ+6ossU+OfbgOjQRHuzzYYl3CPNp
r/vQC3zTm/rOExoPDDC2doq4+j501+DKnKoWgB5JOvBnyifRiMMUMZcgBskf4I4YouSO0iefALrp
GGIm1wf12QDenl8Brz2JedkO0Q//HukH1pIAyNS35P8iLkUczenZ1LjKmaJ3irHsz9gQuivb/l88
ynjI/U40EHPgUjNbpVmRRDh1lLI9WkILBzEMI1K2hMchCQyiCqQ4ahApKQpMq+2qOQqaZq/Y63Nw
cq/Y3dQivLgnWbPEQxWUe3qgvoKAJag62vEhEpcrmQrH8bhvj4MQ4RwgqtfPixjj78pv37vPQjl0
LwBKAtoKmmGVPPZeMiGU8eY/ECs0fktBhp/O/WJ22SYHGTGrUkRSqcE++gRxmz1rC+bkpJN4K5T+
wQDEbzFp7NK9JmFFfZAp/9T28FRysg4TQllIjIl95I5okeLuPZVjCch+NMSf4vdhFclkc598P6tU
ri6S7+IZOONDzgGTLnoY9fR1PD3WSCug/MHx2GZUXuJ55oDMjGAQ+NyUxsvNOs4YM3XkKMuG9iZe
iG6sCcy9tZqB7PPj26fZeECmw/hofm96S3n1rjIwlKuksPtglCtTK5EFxcfZsZGRTFC6SZF5jSdT
gk4y39jIlYGYzVxkvdwBjf0loZaSKqsbP8CWUxfDKQ9HxveUdUF0nwGciy3KBKzZPgBbJKwlsUkA
An9NSLhHUgNA3IIyO+7iUO2srEqO9QPjl0SkJWBUuGegXCJiCbiWVprThyLCvpPHtP+EVfu8E4N1
536aa3K118eFALGpn6FO7ishYXth8JF2rhjcgDI4sA3+BUa/ChVa+C8iVI3wdeoc3RSGqzmQNqHF
OKKEGdKKjyWpLyktm5cesuSILvLcjrtHLlLAzbFSB8rBZHffDh8f5Z3HBAXxL7vPyPD/AUqVoAB0
m9pg7Q+uKTw88mO+ij/CdjJfkC9s/GcZ1KXspTbL0WcMTG1+q4TLzt8aU6OWfg0QUoEPvSv7HznU
RewU9TcvPflXLr1SnzA5U4O47rXIvLzViS9Z9EbJzDUlUqVBXaUE04rb5NSl1vJLiVuAylTPsDtW
6J61E99zzbmw8b/dvRkJs7DXH4OUaa1L5RDZ5UHO3g+dflETdnW3kHjNKmzPcDNEQww3H3VWMRR9
oln5rmP4C8HFSCt+ipyihd2B/mXPHq97uI1jR1W4MZtsilsCK96B5Qn3rpDghPI20IHbAOPCQPGS
3GdtkbNZIc57YquRd5Zgdq5OQFqRGHj0savoZZuydq99kDLVm8VayqwgEj2YxZdqzYmX+zrcRJMv
QrUXhhSjkuUPngYiQetLOS5TRquTyPnZzWjyChIPpWQYY85S23gqLDV5XDt9aA2F54bv/2afTDSX
JwxJKnejShgvghr25nIhviaiazy1KN8UJK5/OwA2saHWcHnk+ySjjaIhwin5+C9vzOsz4AXz2Bbr
nTlX5c3Fnj6OSZhrd7fqlVbzZ+kYQY1BMSJe2oOhHTGf0KIxSpGMgQeiFX+3m4YX44jAelsx6pfv
y5eG1blH/pkYpeoZuET2J4YoPoTih5BvHJUBN+lNWGjGBzSdUTxiDx3iyYnX3pgw371srmRajZX7
U5y8azH/uW6+J1n3bdNgEn1dBg1sDeFBcUnEQLazJ45y9NFtsVNcuuNuHTh9XjQXP7FtztsSxUKO
384Aa4nakvBRPbf6cB5RU+Ls9R5MESHwIuomsqBwB+zPlcKETEC2XxfIZpri8zSnXEi6+Fz7wVOh
dOVMOZxNGMNZxA3t+s4w3NDc1ws/Bip7WdIU0lp3W/rMoEO0hYPywzzmfP7E7fbxPRQcct4F6vk/
2WweOxPENUkh2CWNEmec9iFidda5d1FPiS8qL/U3M3alxSOSrVhHKw8K8fXBkyjl+xRUZbzxd8St
o30G8Vl9IabPodre7KtsacJdhzc+aWZMXSRknHYZJmr4kTUEkiJHimb9dAxtoV+zhjwxb0vYPcqZ
8xbTLdCXJzPwkPJKsFdNopvheJ3gMxG92xSecRy1cQs4PCVQnnP9foDqj5WX2McdJ9MmMPzQlYhj
Z1q/AKiR73MPrzb56GxPeZNPfCxXBihz1qf/OhVdSBQgYYc20/SweeGr5BJGzC6sC6uROcMeUiv9
aK7+Xi6IFdshdlr156JWOm3oXkpQJMPL87DkZ0s37A6BdClnbibMXAF4NeRfCfBdYB1cnzWIheUG
dWHlj2QpDFU0txmAfoZQLrNd+qUQpi4jPxKhjLGnV7AIKKN4vXgR2iOGQMF6UIIvA+Hw3lJ0D7yV
KOc9o+W2qX0Hn9h/+NG/UQLR1Ba5RSzcIQNA9n2pt94SuT2K1itvcRGYopEXW/f/zyxu5Inl/2xc
OV8qH2UIgWBj/ugLJj3rw19ukfaPeNprs/YkOiRFNWpglwt/FQz/sdoU1UAa1QZeCd4uhCde2SJ+
cvGAmeteClWob8axMVB/f3X+4DIgK20sMYH/CdEhFSxlWPXYoMhhmrogi+ioZqFYPuaA9fCrSCF6
aM5Vmp6u0yMNRk8PWIwycvpNWmEVGBxDz3F1ZKTgXE0Uh48YhfNG/lEQ9Gf/o3weIBm0wsiKNz9b
o4j7ctPU8oQn5kYRI6l8fCjlk8oCc7R8spjN9F8OP9JSgJrc1uvhrRODJEPVDleOX4mRfCR1bPXF
ziqVc5Bo/zyglY7y6PqAaHqbCix9NrIMSpWkljSV6ATv1uMiwm7lVkquxhXxA0GZLzqO33X/jKBY
L3L8oYuSIpqZ+RyhEyqh7cqdHwBT4eMmFM92FNBf2DyuN5ACb3AbbkgDgtjSEsbzhdUEP19azvwZ
PBd8aNfBzIdAugsQ+O5eKDkrJqKSMXVEAqPpg3WByqUUeO/4m4VxASvZbFJUNWVrSjr76G/C0eFJ
T+6iXqHUq2W2OrGFVps2MW4rGpLapkgxnOPlZqZ5v7TUdBL1RNWu4169HedtX12TqqRuizsiwz1G
wcwNhTTS9Ixj01pmaIfn4lAbFmSxLJK0y15KMzinPYqRMKXgCzNOyfl4ztwvT+p16FFQa088ArnZ
6881/AtD/ipeIr2VeznHq5P/YSoC/Bmfn9l4A5a3kwXsbw2OtNLGj0OLOC9ntSdRORyb6aRvDno6
tJRx2CzE6OsrnHPmxHK4gBDKmwwvIygV29GurYU79WhACvi6yq83CdGvdP/KQSes0PIvrmBj0/MO
KOTcjy0VSqmuS/ldAvN+CwFsajIkQSX89BLxXNSSd5OJs7rab4dQ29fa6PAgHBPgyK6EnUV/PYLK
UG2+c4SvH2r+eJqVlbYReayKJ7C+Dgd7GtBCENVEppaFFsxyUIQg647D3etBySgEbHcohYisyfPR
5LL8LGBrS4aemzJB5GkN85DdAVq+0JT9Go1XzExTSRK90e2DxkpjsfeQ3bSaN7Yq8zXV536KXZNq
nVnJ8xGFBBixdu4FOqdVD2mt7J9uthHsdc/hYY7gm3JlPnXxF7OQQvYYvJmhEeWgcg9UaQUB1yv+
kJdJvECO7P6TdZ1ndSfxBdwtty4Mq2DdRc+HCrXrfxldaIimcaHHceep3mimKYM/fA1US9UO9yu1
gOZP2Y3Ko5PJliA+5BkNpHDtmHcx6o+XxDOGsZ5nzUtH8mJQkHCK1uxV9Hw57TQtjvxopVDLmAZF
8UFTIeOrjeeCuA9NKj0AqzgvKJfmF3ViXS9Kk13WefdTfgXZ8VpgF7UVxI9zB98XnktwoyfbXXzx
irmeSKZxZ0kD5/OstxyL84Kw7B8o9TjxYTYSFuDmy6F1uv6kQqWB6C68DmBzz58+40usbqTawLyW
/t95Ibn7pKaxZiqazK1ckE4B4t0Gpwae5Gsf/QAvh4alaxxPb8KPKGuRG13e7AxRzv3IBxcezLqA
wQJ+OS3/1z+s8m+6YnqQnOoNorQ363XgLusthMDDCLAeyHFgNzj0ZAYSICSIQX1ovTmsoJBQ5lKR
YqLwRg82EFnQDW5kpULQTr4+PPbQ3FJkY2dpcFINvsroXZXqyLPh5EkxcMRwqkkGjb4EFbMumYVU
MLRdB7TnicPR7OGU6Ybk9xBgg+AynUp2vzdZl11M2PKNfESLWiEuxdQ3Ff9tBB96FyRAMCKCSKWd
cSXDwdKYvqxv5MmD9Z3q51mLKAPL0jw4SZCVgZmRqLZWcpjFp84rbLOPIqs5wOCf4HFVtHZvMM7i
cN6NVCeIGeHDUWIj8CR8EVbhHUxAnDzd2IoFTyTaw6tH3SV/0keuK5QlMfvhn5lWfGibbhkueArs
LixtiPC0WTR06FDmxFuM/pKTV/FqiQge1PKsgcudKNOogTPL6sZXUOJIzbVYcjazIabF/5D4FPlf
7GwdUdpEKDnsDdjcQw5CXs8I1HN2sNLnxMlw7GqvAGtUMB4RpqsEBAx+cTtZdkKDW6Xg6pMnUdUj
y1N4SevzXAZ+D1QsbPLYUuIeHSVfEosFdb6dOKnv/QDPu4odqPRU9iifxVI0PzxpF0z1aDlNspab
DW3MLSCZgakjbsbBjf4NGMFW08rfnh8VvImPDTn/wUAO6L1gR4SnJoP2k5bdRKT2PZSWV+34ORZ4
3eSlQ42wYDVRCyrm/Kx1IcvKgcCYzLpI7c7gHODw3arHv1TvexuvXTjo6bHrivxz8Ke0XT1YOdGo
gC4VlWLrWt8pd0gEwbwq8X0S8iELdKgcw3lElxLuBehdsRcV/Dv77dLf2xaNCtGXiuf8LQJj7mYM
AevOlX3Ab4aDM6cF3vK2MGm72tLarENQJ2RGspElG+O2M9G/S0KtH3jMVSRJ3VU8uWNgx0yCib0p
MNuHVKA/5c24QIv3Zq4+k5biX46rtfoCzHmFVTWHzExBTiMnKdwcKc2uGYC81Ghb4GTuvgI/o7aO
vCotFFvB8laMNyuoXClseF/A9ee2WLdO9M+9efLYZGshdfVO7uwTQCNzDFVQ0yO86htQmkyztCW/
CJKd2dUnFw/pDVAlBHTVwAiVx4kVcO5VrHXNCcIwmWLrUp67jMG0T75gsbb6LG7OU4ye/Br1joUR
yicezHWlCdMMuaMVP252zcltj1G77wxvdn9uBdvTRMrB1wdfWGhrR2ISJofNsFP4SxmYv+O5KU3l
jSaMBLES3PSjXZ9JMveAnGJmZ0CFCx/nScXJfCyfYiC3GLabSExG6L0uJl2VRmZKmcW95UwPbBvM
q20gNuIGYmcc+0ue5lMt7pNIHF/DYb4CwESyzMnzbT+h4LDLXWPCJOg1uDBEp5w93lVjAsYjZoj2
ONJAXrCnIQzlfS8CY/2Fk22mH7ZLrJniLX1kTzJcOuyBUnG40ZhwtOko/wu0HRgQp6m2A79NR49f
d0lT6QN4ooXWCaLmPKRDidi/NMe2K28sHLiqouCgehtVjt1G1HkZlnOgWJGZacToYGb9bxKS+REX
6DV03gcBi4gSppFIPXf8HLy9O8J7fJ08+fZjq84a0wOf2mZRYCnBFdmk+TW26LfO2WM3QhvjxT5y
TLdM88XYVBI3B89ELwUFE5wASDDh2/kvdu5QmBa3C4ptsJ6espKP03DRfq36wmJyKyuaDUOFHzXV
qXk9Rut5Nv+In3/Zvf4IAMIKwfvM9QhFIIoueUPqMY4usbQyqWdxae8sfCVApOUbrOtQwxmJAl+U
i/a+aJ4meTOb/+rPcTQV0Q2zWHVyQhBvMmwuOPex+oT0ZGUSX7/7eE7nUMvEg2R3ih6sRi+ehUOc
T1l/NWEM7HI0ppBtT/jaKm3RZg6qbDqJPg4e5jhBodM/o8H1Pucs2f/k2738jq9a/gNxqOgdRjhQ
+TJ6bCI1MjFytSl8VfvT6cm/vZx8eDrR+swuAZ2KCHer5Z1YXS7c/zJ0ijFVYAq2vY/hLBLRdFir
g7gTNpe7exaNYnqZGYi4QY9eiKwxWaPPzSSqVL8ACUTlv49B1LuHCgh6z1eRXayKGMhlHVni9kn8
W81pY0pxV4jGswK/ljcIpL0lxYGqmbubqfhaQUpCEAIV5PGMWcGLNqR0i5+T3ea8WNuv9BF9FE34
imhKAJ8kJZhcDT2kqfsvHq7tnmIf0XJ34l3MRQYtPiTEjd9mUlSq5WzgJBwmS9Ec156ihx/2LBTO
fCvHVAHczfH9Ga1UF5XW/362gbfQLS0GdW+C/ooxiLMSSVpn50gpipNCQ/vtK0ivGJfzKeFPjyLZ
lkgOPIEWtEfjc1GBsHgrPRF0DhL89ckjBqWjDsc/hq8Mdlh8nutkNzfmgmKrxk8Tfc447XxfV5dU
9luCnTHiLwS/gNmiWXVMd+AK5BW/G1ekYRswB9sLG0+V1U7n6RudBwgU/6L58lZ+LvgwrBis0qWW
Tvtyu5B//JF5Ljbqq6ERLrRXPz0KqroON2yKbNHRZ2ewvNe7ht4TPkXyPFjHXAmH8x7A7qCpynSp
Jrgd3daIxi7cw+6kUUPYt1w+jGCY1mmqutjq9LSehnqBYyDD8YPjs4dhCH1uuZ9a9MI14yfuhY2A
PX88BSFIofjr1sCF8HehIIsyeNStvECA3LZKMMuxooY0QFG0P2QIz4n3mbGIiQPJPMoZ3kIOgxDz
6jHbpu2v2LV3Pi1tUVMP3vlvOcn2DHKe5Jza78rJb4NjzKnocH3KoznLNVvvn/wOlkidzVYdyUoU
e9WhEbslkBaU6rVZ6KXByBQThu2ksGli7z0H8UshVTl5SdubuMpid247PHTZZJ7VwoFNR3U0BpY0
6SrCFfR/LjB/NoqqLvyodexBsMoLrQTN65amycz22S1A8QpYgblmrrgsvGBNMnZLo9RMaUIh3yyc
+ma3K+eLwTA+SdlD/+77GK0j48BfTr4OOXLwL262pPr8lDS1D5w3omCMnI01up4Q+lsNtA05ELIi
vdPenbjYNB06whFizxhbq3sN1LnL5RQz0nss1KVcqAXug7lwASo/3/3aJstkFLS4OdVLfd9aeY45
wrYnBQkjZs83W8doktQ1Lc6YrChIsUUrt30l9EYpnODApdD7b101yhqUUd8oFFk1G8sbn2pnTfWI
LUZhKOTCRHeMb4bV07XNLKOHTnYQv1Wkihg4KOYDwBqmrxiAoT6pNlVJcfhmeV/v5oTfkc0V1ATj
1gGSYGVz+4isXNVbcewIhV2ajpAYCNRtXJ4FcVML4GGFk6f8yB1hrr/k2Zew1PjQ2v2MFQYdI76d
bR7AqbGPVKGu6vTF4fYTW9YHTKQXnZat3rBAJLunW/lxDpcELeu4mVQ1nLOQcrWeMrdro/E2obMO
Ld4lqcPAQF+XBddSykqSK09zaQZ2vAsv1UHEzsWzWQreuTIxBqGzm6Hkcpa6PMraQTf2wsgQyKbG
JLISg8yowPJDkC+jUk1u3QsV34i+aF21xeARE+j4Ke8cc0MraPDoQwrCGVdtYa0cpdCYX/IoFig0
cgqr9XPQx9WgDCoT+MMPaC5crtmvq2OTp1x6nWjT/f6NJlThSswV39Je4f0xDFHYwzZFahST70Sj
tNTWHEMUhELpg9Og5nomqXcv7BfxFL141b90mk19QjCRTAd2LOjLSiAuFp6pJ4HOa/zcO13fQw3M
6GHdE/OeCzNVF6V7VqZmVsurwGJRhhtNc8Ui8CEO+OJrlZ1tbzVQhfXQE4k3kVmVjKdNL5SYzoDd
M/yLfuVq/dBBEf1hLzs1fVol4fnB4Leryl9bPRP88e8+KB1oLK74fDbOWbmemzo0vsQBkUj2e6dR
TobBbzqBg0DVCIxBQWd/wqltr/tjie/on2/6U4aql3l5izqJfhc4nPdaHcnBxrTqVPyeKS+U9Y0H
B040T627+UsobSzxzXLrSBb8Y71Vw38Db+OrfQwbRzelZphYv0OqW6WW+bxTzcS35TGI2L+Vtrvf
ZosDjRTBS4FBaGbMyHGYFg1aDrdyXIQ6BSyaa4isU71RIS365wD2gg6Ts2b9kFfxVQi1nM72C+ze
Tm6muVGSVbk2lzow3498uRGzRaqnbMP1wmshINgbifxoonFG9zsXyvKJnspqp+1fn2rk1upQFc16
zl+g76c9Wsax2keQmG6EoL5iqJp7tXtdCggK+6x1e9Y+hBKBVdTFG1FxCeTe5KnN0w4fP5OgppHD
Zo/iiPdjcmeHk/uwls1YsFSTBDFmshstDXt/TAFej1GrY30RjP/FGtE/I9zkLsHZ7STiOgJzcwL4
Qr8V17k86zw7z3sjJQwt08XVRBHDAvCe9uYph5Sr/AHV8bZaU18M3gkxxygNSAJ7hLUozqRL0th1
DpsS0GC+mcioKhLVGeXbB2j7hR3yYr716DZ/RTifh+L4ih+LX4RW8Ao1Ci1ZQ+nQlJ0N0pRMWyua
CO1yJ0shfgz7d2QEBRWx9lC2jtOn5+GJLEUuFgNAzeTfW3/BmbtkWVzKbfPK1reqQ5+LN5k2pcPL
Ql6p8FELhEVBxkADBcij7SNZlXJ0cYuoNyrk8JuvteT3TWBJxDH+UFu0UOj34jmZJG9Ezw8ztBkK
Jo+yNKtbb4DyAIDE/gSYGqLpMKm5r5mxt/ih8tpmc6x58znxSir8fRnfmoxCqTfzKqR0imsTNrR2
20Hk0bMqClkdPsHRakVZdmJgqfi7key/Ds4KyIu07JI+JZfy09HWqRL5rMOlK/k4Odubq8twIiBV
jIBy7SGPBlIYq7crln1aXqN/LGO/BBRyhwbdBXo5nc5hWKrl0VI655yibmlNF9lJuGFAksdPonKI
R8jPdgkCc+vLRorg6NEVCIWhvXRkDRcXphooifTsv9xFqDtgAdmBiuTDstrifHEYLgrKIpHSQbcl
cQ+eIc5E/77jIYAVnJQkIEMblHM381TnVqQQxWHBDFZFDINEQe9k+suXZmqf0bDqjgDBzidbHBzT
ZHrp5nKpqDWV8IiJfyRDf3PPh9aXtsJZ/wDn3UlynNy728gB+AZjLnAj4sqiY9zAT9dRZICsG+Hy
dfapFAkMbNNwZt0QRtsdnuWEHJ9I5v53kxypMRGkNrSpaOYEzAFVw9xj6Fwv+leneFxvtpsujFYL
/DP8HKFV9TgvNU74HnAVJpFckmu1I3etKyhZ9MRqz5vxNgmtQDIZp/n57F5rMSJJdx1zucCV3opY
BooJjF+6MAUTeg59+PRoif0LqyM61PChSEhfmf/yn/TXQB4C8yN7Fltc8YLV/4d3cPauK2CObdKk
7Wa1nQ6wRrvomMob5aeR0A8ghg+Psjt3bwvsa6YNWlTtQblq6HJvFHf3r4Kvgi2guw1o8Wk0dW8O
Khq7Jxj03HxfI77duDPpTfexgO6tTkqt2Ur9buQL5Cccf5tfCx02ekKWt7pnWdoC4wd8hI5958Lb
uFexLuyh9TJawSkN+ILQ9Vz1lY2gG1hHk41w+sPCyt71rKls3hzkfAFTGZDbHikPS5jb7bQMfZKB
NaaZWJKJOpGAaWPf6PjHbb2ZjgRYe2M+MgKJE9rZjdFDdMaMHckcoYzZj5rcf2MVgu3cU56NRDHf
J8m3/QqQxC7ZhciFOAx/jykALp4EgIyWK03DK46t7UX3XlaeD3dW3nvvbT9+XwBV7gX/KrRA/NSW
Xa9g9OmP6s+tYf6qTUSDfcL/ang7AOtRbFA/C+5R63gzy20DkWr4j5oknVwd+1cLuw8520evhUJ7
A7cT1tnDMqJzitvFdknlzpGa16iJHo4rPsV8Qz1FZt8DYdOeCbKuHKmw0itwHusgaOCEWw0CoUib
9quYrSlPIFLSjV8djk0WSa7laXfAzlYl5tsZXpReET9L41XNrfsPZhzNlUFba2dhwwZCwb7rdKrJ
3jjFgpZoKN/FCmm6i3kyCuXTmrF0qxAFJhYqH7k0XU1kFxFT6260ryv5GTKqE2UJhtIO/3r7S2sV
PGS7i4JW7dcRzoB7J2/ovPErS14/ntp8pPjWKWb+fdDZLwvXtPt/HweAHqTkvLAx8cIZisv0FVSw
Z9cQrS704A6SyNQtfC/hxGEniOYICafV2tihpNcjyA2Xohi2d/IU6sDXs4M/4xItdznsFHUeCPkW
UqNZHYlHxKNlhfbY3A/zmIRpXJuq5T3Uxzgypcjt9/RtE+uIdhAINEm63DieRshSYPjuXfM8izbZ
daIzO9JpVR1oxOU0RqpPvrEbths3NbBRUJrUyt+kplLjKY7RXAx3EjI9FrxPR0M8yWAmxV6TQLud
YZY1dWuYtaDS4aq06uuTjw1xTKV9B276IyQWSSkcpImarSgElqY0JmSzk0mnYvavBRQ+gkrPp8Zg
lv7DTZxOVqTX+gYlfN5C5jdgbddszKna5BhnbLtXtZH59pwv3Ywurj79xuKtOEufnieYGFaE5jhx
j+YaR1ieu5bxWUZcC1HzQ7n412VgMi3myycGKIIgOR3DNMz+3PicWh19v/SriETbp0V3F8Uu9I4f
2JWxLmqCv0xHcPWBFwYh8vcPGyzz+0lIDxADfM0WHmEs2gAhq9M9rdUGsLiujJDdaOraXO87cEaK
ofHzDBiij4NS5oiaDX4+wvLILZwD10SZWi6SMoV6OG1/zk62XNIlSFr845vlHoPfc/V8Vy2p+lnf
TiReQBwgAnE8yc27joM0baLi++IqaNiLgYtPeC2MKIe6Hbwz3keY7KrRsm4iSLD3LJfqGoNYtRxb
C/SqoB1WS8pkXZ+VlkSG4zpMD3y5YZaMSflNbq00zKrJBr5nbZr0bAJlW+lVVhON2IHhomb4VfLM
T9Kc5WzJgyw6Ec/dyQKyZ0D6CAUJCwHuxBLhcSwsDyR9SJrC+NvvXWe5tE4x1Mw3BbKF/Y0YrMYL
Po1h0pzsJj52meDm+YfWMxKp0O+ABiVtxz94bUp7lIlrsaXIe49QUYFh5i80gJhrEaXSXECS9lhv
GdcFZLp4m7Wg8tNNMKOu0JO2/JN5PfrbxBSPszXCnJNDjJ4KyeQadfl6CNyqn6iVjIoSoNe9rY91
z9mKcJowB1y1oJtQX75tRY3Kr2k4hsQmEhyAGyFwN+P7aO4zxXFX/BEyoMbldJnvkZD/3OD2iE+k
hme5qxz1LYoGlzTKvLgstxdYiIGasi98XdGgj1r5XeaJyaE4WqfxY9p/UkJ9f3i4Zb+Gl8/Y87q/
x+iC9jIL9cYB0DyJZpQqON8/qKWbv9dQPfVw3gFdlPQ2vD8RzM3YO/uOCC/UHuZljXtpBiA23T+X
EKREFVRCjvhyGkkVabXUa1gXfLpn8MDmdTbCnBONo3u1bw/ghJ/SdOpHqdMHdGRmv8XBgd7qrJkn
ltJYmJUYZz2XaHXym3q7+ZG2u+ZqH/ATHIHE3dwQLa01tcWjWTTV7MDEMEbGaiV6N263Xd5kd9ep
oeckRBKDraL6MHh3kqyk/DzFEVWxSdMGJDkXjWjU6biTDEMrcIkv5/7zFTt8qKVRf2D8nX9/UZ+t
XcL8MixmuaFk9MRCPUbajy1ZO4ooE4FYj6dtIzeOkCPsif7U262ydOnfc+SNqB1fLT/VkaQYVAO6
KwADqYHsN4Bz0NawRdTQ8Qzihq+VLvmEZH7v6BEXJ/sSbAiwqXrV++OLs/7G42D6NAxuf0MYRf2e
6mhG83vZ6imKqthOyTF/v6HO48bDUEjI1s7h08Krh5Tusb/K7GNylRqxNC58BCot7tNr6D5LCfAW
RQjj/MwcxSQH0/5appE7h/nLDDzEaD1htKxWhieof9aBtX8t2GzsAExOyivHcwkwsLZjXAWE/ZAs
NiM5f5OQGAGZUVQBNmSGEPUO6JbKxPzv0MHyGr4yvYutJn5jZ2rq0ZtITY53MLfkLqe77rjRP23I
RXwtIkUMHF4Sh+lK2vo4o/awkaHuN1Xn/Pp6zdddBuu8Kc2eSgh7fIxmbJVSlWewyOWmgTfkth9e
FG4dG06iYYAv7BGTl8ncMIy9DQQsViA8S51GW5eaGOi2aBCVyL5FcUA9ZlO4mRsyXRpwXiiS2B3J
WVEvpdmS+ROgRfAHOOyuES+cxtYwy0++T977JYq0w/H0HuQTGTwQRa+4sGpRkoi/klbasW/XoFHr
cZR1tfvdNvz17JDyrZEjC+2qB4dcT4bJDc9Wc6i9c93boBPiBA4L7eJaz0Z0N5VnCdMWZbebNG0E
rYW/QCqqjNXYGvj043TJNftaftzGymPCQYP/tFxS9VPQZEUZAZ6SDwbiAazqUewSz/x67CZyaTl+
oZWXM7toi8Nk2kI3CSl6DDavzHZLVFEI9clCUEmpThoP7Oqoz4J73p470uDadzTNqzdxP24n8cKw
DiVbNEG652xzVve5wpZHMFgFy1Q/Lbh8+m2jmgBTxQItmaB8wMahSHFqP7OHX8WanYVjmn9pcvfJ
z7qaiOKX6ouafcilMyHITWnjjCPDXbbahKurzR2i22hJBVqDFI7FAtyZyMh12ugskpL5o0/u/kgY
J6GRkftXf/XwAhjoD7dEEQ/+VQlCr1uOespNo+3l1wblsgGVzzfzwo6FdRhx4qHgb3vvkA2QItaf
QkAM/kh0pg9Os2coGgD2JkrqfcOt6q/Hxfmoyv77fSK3g1Th5p6NJvLPpP21LmRl6zUM1kA726yV
5B9bf6c5i5Dncww2Oi2u0X6WPwtmXZQKxddlfCqSTRN6sbYStVyfi2fabrtSbn01eT2MB6aN3qee
jnqDrtD4sQB82hCKuk2OYt+15A8/uzG3Vay/0S5rz83BifV5sFcYDCbEp6RjX9+brbBVsANYUksv
Te1tIqNU11nYCEehbYTBLDijyzM02QqcYKIaaUgbfBxaBeLaiUqccSNYMWFUihDxArykxYc3kJGi
fnDnz2CwAXCSyzENu8w3QVT7E3E7nlYD/1AVGpBEELjPYdI4Sy1r+p0RZdjC2O6e7dvMwboNS3/y
CdrB36i1/GVtj073Yh/K8kBdSp4k4OGMMJQVXCKOGwHSafP1vyZfHBoOoGG2oZx3ZfVQuUZS99YD
+hbGtmVcZaCDcskeMI2LS2nl9PvRwcTIyHwY+nXGmz2nAOA7ou1FKtzfoj3i7V2qdTYtOkXPucER
+lylYSjtCyQZXP+ajbh/MnMVPYegJEo+XDA2UMITxH0dNYRfjXdnrjIZgfBizagrGcWJe+iYYHhy
0NiuSL0CGX/geAsby+ysXE6ZalaXglMrZ3NPwymP+fWSnBsmmQkTI4txAVH1CFyvqSSjy65AqWY+
JAwRx89ZEvqajaf8+rkEJDeKYw+LXqvtdEJxaXCew1XhMLm1jwFK9INvPOSzVX83wNqE6FGl5oZz
GgbFQM/9VY0GqQWWvjN8vRyh4QkhpUAcr8Zj0ezUzk4qMceaHwue3tw/vsR0dM5nBViv57FcaNUV
cL6UljEU6TKcAFkLcrmR4QK17V3Arq6fytc0lFkbjP9ITj7oGMGIgkwrDE+3hP4b0kCIiDqBsP7Q
ClrM5Y7mTOCw1wEzcRkC0F5K6Cr9CKCHkIAXK2bY1d1+RJH2HY7lW9+Khu/I8CLn0TrXs6t7ywTc
+V1vFITFrpO3eTkaflTrUdf+0MxCU+prBonSMNUCCsQWDSm1eKfLmWN/N4V46qciqX/9sRABRWjN
f8FYw6XaDA8FWA4Vai78+bobew+T4gtfUgY6y02/B9/iMLtjQnyXgJiOK9pOymHafJ3dDm0ATd+T
F3QUXXyPPAQ/mF3WoFm8Hfn8wLMr1YulbGpSF4J8MoCz4nHWcR17da+5L9gsgb2PTRAKW7Va9OFn
P5mJma25DPuKhm2SbcsV6fZIvvgUiimG9RjIwB/K/e52DV/NECVVHvdglgAXxrg7hWaXIjgccYBk
96ZDZrteXCilDmMUoPI+qe7ue9nwep42mOtiYOs4Yse5UYzLnTmQA7toWwDx8kuy1bHv+z/FOFD4
dgL4OcpY1QlfHrln1L1dBIJSOXS+rmRvap2ONvJE2bpN0XpfQoEJ01LLIn+qdz36VNpKbZuaI9s7
YMcK0OzakAw4JRsB7HCeGD4nf0Zap0FWHogYV9nRuVOmAfeB0N3IMFePKZU4zWZTa/OPZFcBTcQg
+PWpW6ueRgeI3AuWm3WP15ooDZYtH6fGIoZOoEChBz3kq7HnwP3Fk7/WIYwPAcqJ7ZER3ufbIxEr
9wF0OzfcZiTve3s2IuXNRysJDxpYuQjfTO7epouf5iaVk8SksspGO8My6GXC/FaManQWF2uMquPF
i1exBwFgv5t11H511o7ra7rInkiJW8qgJ76x3YAnVW+Ilqw3Z0qA039vD8+ZMCt9ZkBVaxDZAKCm
CCwFiYItz8kRN6DbBU2gC5mo6C1TRyUJeix0zpOfj7Uasc1BY3zzSkAVT3zqryyB3xunSqHptELt
a68CeUZ0SNIT82hat00u+SAPWLVVeuMyFFePoI5baJM8g8DszttLfRCoKlKxh8GD+aG/WZ+Q97vO
zi3Os0CJ2PhJs4OZht+xW6BSYxpxM68kZO2T4PMV2lclpLymRDUmLH6COBr5wg8RfQZxoMn+0DuJ
oHSGrd1tG8XMoHNejgfHODbUIlkn48P98m5ILSpCmHcKKQ8PeqwdVK9I09LGvWTT4URtGxx+ZkRc
h5bDfjHKAJzBJ9WpbnXnQGmDj9NmSmin2dkmavb9Wbr2njW2KM2fXabkVEkdEYalgCOoXUlr/bX/
orNbIvfcTjVFL03aS/fajwHqr9qryFhF3QZnBVB9Q65K4fw2/XTarRnQqnBVtzydSBI5+qvQPGz6
3Ed/EeHf967DqC9gYu5Ay7sivvhjIjCseZT69FsyeArK1ZqYDvw677HehcY13vWTX+Me7a4O9A8q
qAwXBiEa9Eh/XXuScHqRsu67XNrzTCd6NaJJ2jtvQiIQQV+x9K5HUPukJg1reArDcCKcRDPgn+qY
gArJjoePbmuXc6O64XkSEZx/fgZTK1LW4zdHasmn7XPxOeNaibY/K1DaFMwix4PkDOZwpi1R3Qzr
s7/38++Y54QPT8OGxbh9OMwB2nnnRN2oaglNc4ZLzEitWMsX+c4/REbAUQ+RBgN0KsySvaCo8evW
V1WHE4TnE0a0LPVT5/XMkCEjBCJrB5PUDjUMjhCjQ0PK0mN+XhNMw7BNSPU93Yw/lfmaJsIM//hB
PFvHB/yzw1TwlDrtbNVhFycVoThBFmkdSFM0Jl9dtN+sFEqusM/7xQTFYC1XpNoCLkjuvqu9qEsp
7FyPqJ0Qlt96u9V4m8x6tJLJ7N79Ga44P5pw49y7/heV0xrn/QFbTPvs0sqPmSgc7yZszryqeNyH
2M33YnekU/kqGPgkyonBm+3r1wNi4j+7IYyYOl9o5gg11nfgaK6apmSkB35I7yu27wpyTAPXeTLr
nUNPH+MecwRgRBv23VnT8qs4F5nMLBD5G3CDla5cFNAddFf4R4VBGJkBrZAWqrSA2+ZD1ykQSAPN
cl5RewuSVYDh9Xo3sVo899WQYbFccDZj2Ed/u/Tp5vrhRCdlRiU/OWx4xmk/6/DW5qIaJm5g92ei
ZUuP6DzxTMAAaGrBfJPLyvbs+yJ81Wh5XgolNiJGqtovZSTc7y55fvHXzt09wz7yig1DT1uqaTDk
8fH9OJ9S5/B6Qr4tuT1aNhcmOENXIIX2jKDkIStT+f5AeuYV8o8HcIu97pBvjgiGhoD9IFZxQs5F
7S1tMKuh8xwDiZ4BSve/etDAfnHxhJKbC38eEm1ZewvOQ/7Ypk6E2xpyvAEAxHO0AI9IHcEpmUtI
Sckw5tI8P/PW4nZvBsezl5b7HuXYVrgjG+VGydBjLpbpOXC3ExxfSj9LyYfEdvh6yAzQFZWijXMr
Ylnrllxa9daRFoBqUcxxdNb7x8/VYbx1z7Dam77rGqkjd+hImxcFzZDFfI7Hnga+ldNt8unPne7d
McHxL2B9n0DtuVGLhUgno4utqe8zCIlJ1puVzLsI2MAZlkWqsj1CRhR1lC1DsyWgB9pvWZb/j7vb
i+YGhiBdzI6R78Kwh7ERHMeXcZGa7voR/ukGaVisGu+sdXdLIspjad0s7QVdKqV7m5Gv4seNexSm
1rFX0d6bOMHmYoj77/g3eKqoXyFYyv+rpb0+AOWH4o/bgGDmHhpbcOiqiPyNjC2P11NlEH4PjTME
fodHTIaFZqMD814aOPlmUkHjJkkk1Xnxkj5cm4L2fxZAlw1fplpSZYfiRxDPdgCe6wVqb2FL5XZv
TFWvvoanwakYpUFBdp9gHtYAFq7cRyRTsgoXHvEDhbdeaMFp1c//0jo2/0tUsxMhRTIGtdL53aTl
kdPAQ1cdTYX50mlYn4wh2kq4ag6VQabK6BXO0frMKufsCC7mEejmarIBfiF/9pKqxbj5+lqiDs9n
vjLEp8iDJ8NqcUUWdn69JHDgQwSNFK5ze9Fa18UC+xYxwXK+fBl86AzoPdkCvT6xr+L+z+7+QxhQ
bFscIbWHkLMujEmnIPXBJNqU6SxqxF/+bZ872snEUy25tBr2g2OwWI6R+EWWMW9ArdXc8q0h0OqM
2U/+8vcCSQbCeRQeI6WwOYKLc3LiL5vRvxL/fQcOvR4uGQNqMU1laowgkFbweBJuTdGWg1RVFqiR
L3HCxAJTFzg8B1jlFl/rqaCbtnSKRvyUzTIm4h6KsjLYpW5tX6w4skZeQA3jMqqC0a3B7aAL1Y1K
ys212EGre9vIBoIOgTK1BGIGE27GCpTrw2zpT+3HSQ1r2DHYwcjv4oRAYfa5GSfWMEgul6mBhMWh
ifjNXgKKzxgIPO1h3cnswNUVLwTsIcLpTI75xJr5HMDERdy7tfvxPVkd0Lxx7O25XOAUmO+J8O9d
KSRlHfWN9hQWuXujOdIszyEnxJm9VwfdmBVXrCiKNMBHGs24AVBQvy1KGOaxiwfMKXb0hlWn+rZ+
+SQSRkciEn9zYfp+AkThGExH4XRb6HbovDBQNYTbePkwIjZXefrqIxGXQ2RLZ/rq0QkOJbJrZ22W
ydA/GOc2KB08nBJ80s64v7iTq+FVSUQiktHdKoxM9AgJtrNiGR/jI0r79eGSfMiknbqTkh5q6nFu
gpAZpo0L/RKkpEVRUcaJH0i01vSUYVcxkOGb2BSHq5kKfonnOQLK62bkfgm58OV3j8GInoZyxPq1
M8C5KtgwFM+WcWdlSm3Ob0wLWPfHS1FsX6i7uitvsGZRcC2GXqGbc5cRLGi8PC/ae0trwzxnh0OT
uxVD5iDSWqwmhyvvO3CHYil0c+X+TBd4OgBOYdHW7Yz6B70BSkMKw28TJBxp8thapty7jKiMAOPj
ZP0uVREa/kSNlc0spHW61FTwzSOH6JNu5QCajp0ZzB2YPB7YvSHAvdXA8ew/2cD5oGgdARNxJfFf
Tq9+vay7vGFHz8ywRxZuobjKu0vblAq/OMXfhayHytQoj53dT+QxImNzpaRmKscvopgFeoxBtcvz
PjlBoGVWzoORAFvSl+iaPEnEJQlbpRjM5jEPn7ZsU0RvTojlZrORfF2XdTjCBgLTirkvkDdiU+XD
Q5WTVTeyK+ycYaLIS8psAaPZ6bwgyXP+JDCP2NYjYfrG/SLdjp7Jb7Yg/iEmtpvo82DowHy9JbSC
FE8Z5mAAxr66qyNzs1FwCZqa9WfdET5hT6npu5YaoVBc6/tP14jf1552aI5o8KksTaQkORwSt6C4
Oo6aAR0W9vHmBnGIjIsE+xL8kXusB4j3H/9fZ4GgAopVi3iu3s4XRYeR10U7CJUy9NKRAXXxln/E
wRf+nJ8MPEMkPYhqPNRGg8NwR6NmKs2smxRNF5eZIS7SycelcJBftw22xMqtVMPUKLyo+JlHJkZi
gPvAYyX2Px7PcYvWjRFBpm2v86aypdh7lTCZajFcntbO7zuzc70ir6iz3KUGVkn7gY+hnBUBjKCI
wfREiKrbZIAaikE/Xi0XCBScTMNNC+FxFHV76kuriY26tw7Et4Duwdi8Ezm9EgcPUyHL8dsmqjiB
2HTWg8Ckvj15vdPrZuUwmalOAeE0u7Id+Gv1z5s9k7zXhzNMQ33FkcOdCr1ioABOlEPRalgKUr3b
icuAe+xxN5a5/5mNYn4TWLvHnZTn3+j7KCENuloADLzKmbD6N1jtGO12z8HTLeF7bJy8bIL+gFVM
+KPHJ9hf0dupEN4qNmo7w7EcvLpwXiALMB0NpgEuJq3wBCtw9jeaOBWntrOzdyrlF6jqYJ9tZh/I
sghhOkeQH8vULzvmMyimNM5Fvg78E4Icmh8ogUdgv+0Aedrtvtt7OluCri/EVmbTaXzs7gxiSyBe
Fcr1NCl02/0NW4homZfatjP5IJXL37TXeWAcpMiW5Th1dMNw0facyohAb00vl/jru4XXk/TxBjcw
HW2b2Lr2HK/BH/4aV6bgb5CPjtT4Mqc5XABiSqwVyGT7+shnmiJ1rg8PW5HWTEhoOX0qc/I7aDy9
08eKAamaxNaneEEdY2at+k8BsF1lmfBP7l7TRbkBDBZ16UNxZflQlyd0iUf3RcPc2X5vXnuo+2CM
0VVai0KZnQv09xx8jJrizJ93gZTOauTK5/pRWkLNRLp4iNIrpy58Zo2Geo6OP+V/IjoMhLmZM0q2
EV5hDhDvXEyHGPYRC5IsekkF16JcSU+fHwWRO/w65F3stUaYuCr8Cucs+mZu2H0+wxXWdRtIqBee
meTtCmMDG/mBjSgy1CTzXhWGYkfF5TVkzQHWHqFJzgXytSpd5Eh7d4EhtzmUKAMLk1kLt4eb9wDI
N3XoARniE+ZH/4ozt/bRRYXx5a1dHUu4dl/doXzcZUJ/1ylJuPehckB7GMIpvzFdbQshosK5llCl
nxFtKWCdD2f0i7PaKmPrYGI/8rdtcG9agJnKR5eKrGfz7I9Q8Jq1fOoIuqub0tghjSDiQxkzXVVL
QI8mSh3wCUmSMNelrXEcrABpgnMvcnFC6H4vUaPj/hC7l3acz1BUeHob854kLJby3ACfTvSJlZYB
hQRMKfDWpCXmrLE27TYsXLjmfi6Ml710rwg1GauKWtP5mZMHVvSk3xggYIMENupvAmB2kWD4jM7p
5J5WkuLy8VTfUl2o0e8DIILSRXKrUqBUAphA76EoplfjHZZW4qlsTbRSV7QcDIEe9KlKk7Nje5Ck
I3Oh74Az9vvuxT19NnGcRkV4DLu9V5g8AenmvypIUijiWgKZDYP8BHwiIA4YqH4vIxOwtEB1ELyF
h6w7z22P/zF4I6G1hreipUiwTjxJlfNuF6U+yeqHSHhhqIE1I3JfjlNwamnp1nrtYh90bGPWaAbK
TdGZcHjvg9+BATAvoc1HZfQvaAf5LZMPl7E4JIEEntdPBq4p+CJVDbBPv2j1p1/H0kqRqEvPE/kn
1Ew7aa7w+P6LA/RAuvLara25bAOOTxSWVuhw7/RzBkuOWt4oXxJU4g/WriadfI+ryEpYHSx/oYJj
hIgsQSzadVt62b4WZ667guOZsNo+iTbpW9rSHsrt7mIBqHxLtEk9AdQsNNt7nuHJwmBSiOFD/T3r
29bdwdnEjFr8FRzv8lHUBpvukhZJtzTtlfPH/qZa8A19Gu/RUS7MD2ZgQ3b9+ckYdailQ/VJp2st
COu/xqAkus1dMf5kQYUM2Y+AvOzMAww75NJiB9wiXbr+DyfwV3xW6CSk3/EzQwevD14ebDkKXDz7
OeX+wiqvxlpV5Q1IpjqFx5+bI6H5uzI7bSANfluQJlNxJdzhglRsuuZGYReq6LD8apG9lAslKg8T
s2RygbDRRREbKUGde/c6hiHd2bG0eCowfziacXLZ9In9xYBeLQM6Xb19EU/kT4YriuBoDUqnWe+p
jYPKkWyjV/1fn+7LB+1Fj22nLj2lekQmn4VVRcn3Ni0OixnxCKBEssHor6ERSYv1eUO+qokudZFa
vSfdrxmRAx1756Svlq6/USKM9y6oKjPO4oA7fwb/o04+iXr1cuAWD1bMAJYAWxD2rskeD4S1i+p7
m/pMynAuK/Kxtt0ZTQqKFZWTTUsIgIJYuO5B1YhF3I020ju6hAd/demJvL8muX3aVciPHXBqaWjV
O7CaKeVcd0nPhJ6BQd0Mwmzni3ave9icaZ4d59RlAl/+Dq84mwEOhIT76Dr93a6U3pVV91DpWuqV
cVTQQt85kT2wH/l9CzFS3DOA6hMXt7egqSeDMZMpCVARZR5m62O0WMCBad54T3mVEBGtdRIX38yu
+xe34g90Mv3nEzBefbvBv/eggS3Up58UOmlVqrER+VmdRKWgfgevUyb9W6UVTySFJf8mopQUwsGg
bgKHsxRKyyvrSpQ4bHoMXsSCfjHYMn72COnOMezfhN9DvtSAtb3tPaLyLHBNVGwce4UIOtR3xQKf
UYaHCRxYhrXUpcuJGHR/rVHmRPr4+DY7DvO3DsjgwTuJsgAgDJX0KfzqOiMxk0WmYt8o57EAdd4J
wXnE0iTXc3MPHbJIQZjGMuVuWlnO/+4RatLbm621ddKcErRKnA4HT8smlaSze+6z6kDQnSUoSPCV
N5WToMYpcn1p8acItmLmnH0/ZeAjGReXp6Jb1+36BEWypHTXM3MNhypJGoqVIMb9y+u7ak4pP9cQ
lwcyRwSNO/9Bp3nY6FZ2gC9ab1qW4HNtWzPXThRJIvwGLZFT3HY07dlQS3L5q3RcGRBHE8QI1ZqA
sn1ZopxKEs+XTRTf3iDc3GtoO/kiL5QqHjG6G1/5hjOxOISiDvrESdHW2jbHjf7No3U4jxvwm5SW
EgPO0CBbgLlCWgVmfXcmfT7lBpVe6fRlNV48mU8Uf5BgmWd4jyB08+3pY9R72oBlVGYbzIZpFoOI
UCmDp/rrXdOY9M7aXU3mAF7JWh5jPiYUeaO09IoUsc1fQ3c4lVUOFrSQ61vnBbsKFPH/RnuXe0SZ
etH/RE+Eig4bK1i6GYhE0+iBExNWLg/hBcuSQDZTABRNhwIdLd5r/iCBfrFF7/s43/d1EA65aE0h
G7RGAxaXqWNGc2fz2OZECA3s0GogsUudIoY+88nX5ctfK1Vr5tHJGSM48v1avPT5seKCmS4kAsgJ
oCle04NaioO4xl7xY1J0Gpn5YWv3LQkvayxFCeqKfLJvVQ9trxHqRmPs8A6A6qD9GLAE0X4sxAtX
tKebLuejcWJiO4Bwypa7P0Ok+m3P9GSPKl6akab/lhZMpSgeWU8fbFwXLq7F1/j0lhVMdyR+dDUS
o1ckN75g0WYuB41djbn2C6qQdyscO1TANvPgWHOVbAMMYkU/LH909RuZjFynB6IKdRTJ5dNA1Lu+
BdDR92IfXy5O29HwFXkwAhgAVSjZBkVA3+C1jOLUPJ9RNdUlUVtg2q+3UkLCYdvSAlmz/RlSUj69
OaBonAVSg4d/ps63TEbp0RnB5cYRVhUdPxgSkXkooDTeibhTWsGX695XatMh+KqzbiTCvzOsx6Gf
pw5UftHdNKMDlUJ3xjg+yNor34+0D9ku42SvB1ArYqCyRXZ93PnN2pR84w/i7Zn7M4MNZeHvRIe+
dMag5SH5KjIrJP+eYZAcCppIjCy4nsvYA9zERO5rg6OfPGvHE6HsyVsRg3nXvyvhoegsOqOYuyJf
ANc+4urfQXtZWHoWxVI1grpYmZTou+c3VhG0IOKOzRJNWYikwTCSJW6+/XwTY8Bm+h1PAvh3pFqJ
nEj7/aMaIauhZDvmkuctQvnpA31vSrVFvpfrUSiC4/vJ+AVDnhrzpfFPxU4Q3oF9lXGndshuwe22
f5jYd69Rqi4X6DtwWFrYHJT3HtAZG9EGRdGVUD03kFsNfOTlqEEUmu0ONt2Qd4L2lhF5kuVJWp8K
2we/nRZQlUHS81zm2IY8y/LzPox84vY4FCWeQVMf8GYJCRdnhGghg5mOLhExQ6EI/GG9uN01QLWu
j814aLzXRefKigZXtMWpwUCKuMj6tnOJ3MeUZAXsFgqsOZ/EL4Fbxk7oM1E0Mhe3H0lIHReMu3wy
ncpw3U/jKzggL7gA1r1knLodKYkvX5Fls+kMSiiBbDDEFZvN/QASqAqsfYHCPn3rTUoZ4hfoFQbP
mE8Jb+vWyNdzaxH4IykK9ZRm71lrzb8qiYJcwfgZeyC1zENDTHtfo9+uigGACYD9zxFJfS6X3E7I
9vHf7UH2LFnWgmRiju0lXsFzZYjFu8qnJAWY9Yaby7goQa+c2j9Gm8Bp4JOUTzL2weKur7LHspIB
0FgkgxLqCY20b1mdQFCd+qEtnWpPevx54M6mfGU4M8dxak/TfiHiJY8kyeSRLnlDjkFS7Y/dJ/+0
m5DBInvCE1WWI3a894z51OeFmgn6pI2thBBGU/djEuykD/IbDt4N6pCKaJWViiDdJUH+Ji8A6ei1
B5Kbe4ecOrU4yvc0noZJ9vNGQmn7Aouc/PNkn2a2cIL5GAbnrLhTvc+pr9zhxAzm6IUo/xoXukxO
hRnQCubgzDDalfKss1edDxtvcm1PnlvNKosZTcM36P5kAN4mzmt/3JQMJFAEcKB5W8IgL9vF9G09
xSBXf0BOnnEE9Nj027WWJ1Fuyc5d4wd/y77OEPnL12hUbac1xjaZsDc2ncixcXXHkJJ+Co5/ss6R
qFDlia0pAOEIMTlujOpcOZx9Cjy2Zzhfo/PycHHFNcIC0WDDI19r6qEN/wg+Un51BeDWzK1GT4eZ
OQY5sWwhLxoBKM5U1SIVmAPEux8gkyrcRTSZMU6IHG4VQzfYDG8LpeIAvLUgEma41HvYKD+CzxZx
ylHTGyQyD5xmbmB0BEMUKOXluiF30++qWt7/S/++6EYKbrx2OvThiIVKgwd/RygzY9QG+CP+fTKJ
7LlmX02MktPlbPTHLWE5Pw/Xe/07bSUz/dtyoUdabLrqkQjW7h8EKYcFjn//quzRxd3vMrMdEUBC
iwLdpaNSsGc4YnQ6PF1ozqXwXxwhgobnIPpRhoDwFbxl/Op/0oddbSKI016EarQzVTP0uZJL3meh
olFZ9T9BX0jf4/5G72PDwyHtH5wwl822CYo4npWzKTPgBhH3EFUXcn5Y/3NuMby/SGh71cXbMg6+
xoOv8OSld5pbaMusXLEyynfzIXXNIdVXfALljM8LDPo3NC75HIJsQ5w1Yj9yRj86UgWcXshbwnSq
K7dFCyP5eZs1D3tcBkvcaRX16WKZUjD6WokgoTPsH6YTSVEvwLnlfCDqn1au+QfTtnf8kUe6unAx
0ek2s5NZQ9IIXzRlE/GXBKqriVXky/VRQq21/XvQCkzN2Q171TLR28swwbADnYigq/mOdubWudf/
4y0nBfrOIsuAi+BmlguVYfz77JDegdgKxLxH4ufwNTn8C+xKwUTUN4hF/E4aKvSYO2L1c5H0Sakn
ueuxcBPyvBu+7+jy7lPjjmeu8LnIMLHLZ1+LCHBCNCQzloA016tNw2vKigxS3PsXBwBD7PQUZXUO
DWE2pyLDtpUhyqvv+b9ragjZhY1cF7RXfl0t3IL0CvnWAw5UtThEpNNgOVnV7Lh80cybgw7+0kY9
ywVY1x1By5LQ2GYehheWTa+3aJLEb2IfOEIeYxEgj/7Tkc3VsOOPcTWUi+pGlBYaNr23ACvw7ra7
nRmKZlBlb8joDquoZdMGYGhLxAUmsR5Rtp9z0zqIjRyTqnvgPtbtxAjoIgdzGScHnPqsy2Zwvw1s
Ki4apq81vLBcG2YHOXlwDpbTZfSUofcbtzKmrCmTrFVJzCbGjOtO79tQbcyvHPMQ25s1YfV++bGq
gvBI0XFwrLYdUPUhVTESHnr7YGtnSK2vOGb7+jWAEDYyym7okiAYziHxhsbk6U+nFSgB01Zor6uy
g6iaGkSVhCiXspi7yauAZBIbg6BKZlCrfe6OC99I9wLjviJBYQ5dELSnZpyJCFL0/W7w9qZHOBFG
TnmqCYE1ijVmamS9oFbg7JY0jiNlxmOnkL6ekvhYrjPtZy1ZuG01uq1VnbtUxZnNY/ZyH8nY/kvq
5ORG7GuFoAJYYYM0PBK5jloxoiAItxHDGXz5stkL7Pd9UwtEmE+xXb9kKojhTUSnlFv4aplXrq0B
J+YxFdMh1V1Lx7ZUYDHoeMLhlilpAN6JUTY9XgG+EEt2r4oyz4Qk4HcVoQCeunqtR8LesQae1x40
SntRFD8+rwvE786WEAkowrq3ha+NpxEANTtLdbQvGA0FtpzqV+RDgM6ozP5zjKumuCGb3tZmhd6n
GJ2Bp1ETByMX7XjS1ymO8TvWuNdZKGjzFBT9p0gIPqBmckl7w1KhFSQEuPzMVKECTp4cziJ5d1xp
n2mzts7XeT7SYfwCuCRcJK2FoxDeXowl6OPvlvriw7EI5syrEwLZ2L7eTp48ieEi1Tv/NzP2/wcb
2gUxwBd2erfru5/IQDYZeR7YFmF0o+Z7JIiZI1JQpP304nrXbjGPSueTmIZhUUZ1bvcvogzs1Bk8
Wb5wOSC9hldOKNhFqIQFcXwHbVrrNlCmBMpclPTnLcOE5yJh+e46OIbqijGqi+NHW5QNH2mcignC
KD5tu6XIbUP9CT7LBmmr5eZVqJ8BhV8hFNGRzpL3GnxwM1oCdrwoYB+GXhcMY52+vvrn7+t2WgPQ
0QwXj4akEps4uEnoJuMZzBkjtJUkG4PaDLHTnvU/pz55pJJTenivuwNX5EFVQ1Ckd2pOfaguhkju
IQWUvOHETHj1gz2XoKxxgDwE6gLNq3KXW+86xRl3KgWiUUlSOoBDVGQzclk4LRMB2GUzzv1CAL8a
OBR0LC1uPdjLjbtIhvb5GKD3avE1SX664UjNPYzKzWsmJMn7aqpixsl1mJZeh+GfA1IiDJOjWsRB
IzdPk5/7wHnBU92ZLnyWEVGdrbOH0I+nFX+Uks/Jao8HtZyBJ8FSkjjC/hAAXxPPYGOiCnjHSngH
02Dc7+4NWCLC5+r2DCQFJFWjicZx/fBO5P87jig9nwBV/aTjs4K+NkGp4Gqxry9R+wwG4STpMpfX
W5WAutWXZl0nOnkbw3gTySs1Lo+IIfQ1cXOU1yVG3QNAH+CYDdooGAxgUWWD77Z9nLCAcg/iG6xK
4qv7b4fu+ImAxiIXoCmLDMg06u0v1kO+RslAj2m1c4GcTeqvGGf3vp1G82DCGytF676Qv0cvrDl4
NXnIT8QgElSrJEliAwBeuZoFh4xr84MPGleET9qm2MzeVVueImyuK0Ok1uZFGUo5jKgfnrnbHtNv
sMbOsvLTPFSimix8q3Etn8uK2YX43pEIh+OAgvJNnat3Dg3KzRoIFwBwff3/C47SN9RpRY/FwevN
4cBHP8F0+GS353Q8fXuDBWqBrBPcVl58ybkrvLz6rusGJQ0kkIR0E5AfSPqSwi/MGfROhAUo6Y8w
ocmJSz1wCA+SEok4FnLk/+Ts/8M81EnYzx3Dknim3QjDbWZNWttrKTdyoMT4DYQmdEudzFf9XkHs
heNiY/+6kDGKupFtpBwzdywFZn2gnZss74RSmJO+uFuszfjmtfIHIfmuDemnOy9OKAWqxoeTGygJ
S/R4mBR/5zvgXwWiSrN4Bh03XyvOd/OsG5NcY9pLkFatIFAWb7DbOHtBCyHT4nYGfOy8Wr2+e3wJ
/rYkNb9bdfmOhlS/SAZwKQiCNiIzVSCmrrxHW+koMfF7/Vax7X2Alt3zoT3v3YjVJWC/B+WCADsD
h6WEdywxgBcRaPo/jDPlX2Fa5rpJnqqXWUo9GAcxXqZLaXkBHJzr91P/Y8MHfuHqkhW4Sj3SCb5i
p6BhQ4bBXaPl+zvnJelO0Ht03lC5CGwid//fFkmuqVt9pBOwJSHgS/FN9NJHhs8MmCkJdk4+MEF4
e+zsvomqc8QMUXsjBChiAs7UeM783gkx4tul8i29bMtOKdUliESSGcEO61oSXSzVeYgR0QJmmgOU
RG7ocyqEicdPDGYs4ZhvVNEAuHuzWbh4t5IacTc4w7qmDMz3SgIlYo/q0A3h2bzk5mCq+cwFMw6P
5Igrz4oG4Jx42wDuv2EK1WBN2zsS0AFdTvwtRAPlq1ljaG6k+HmhleHK1+j1++oVQ5NzNtL7mi3M
RzzIBWYsmueyrY+N0urFHDtd/bawcvF32SKfJMcct5cgvDDPoG2vL32PntK73eGiWbZ1GSBhzHRO
poTuryamVKabYzLftfNSd18lrUXgtVH9PkWaX8ttpu3NmM6jXa8YxiKUaS8KI+W72I/wf9X3O8VP
OjLPcxS9ChDGIYhca0cosG4N7FyqAAUW4woGJXOViASfgV5ELzLnsThUmdaFqtSdx31YeSeWshZb
N7TN2+Gd8RKWpVOFtjANFLjPFn/gFJvWL3kDDG2+cnSkvz3RW9sj4HXQEz5tQ6XHl9MHqiTkpO4z
2yuZ3WQ75BkH4uIOuurD0lihKBQDJfn4dU6/YIM7Sc11V54ywrwEW5kogp9jwGyLbJcU6gOdgF4w
G1k/jMeABMqeR09j4edikr8C1XkoNlDt+tD+4fDhSwj20HGwLdhDHI3MW+lx4Wi7afm/2C/IYays
Oh5j1BU9RJmU8Yn38hM7XDUTanh8XJsNeQqm8Eb+UXCwwtE0v/ypOsoP+vvS3oJ4iS2PAJHuzrtH
/gVTGU/s/lydqprR+FdXSprzIFPqr6eqhPreaBm6fn584FzSs1zbp5LaSK9NkxyfK52DGBzlC8qE
3K1Ko0Qc+CPXDcrNyRI3vvtvjmCKwnBQFYMtV2NQeQjmLlMGbJ10wskfstxRfq5BVujuTnK1UJIq
EFymQdsNH8Ta32J7Q+9XyRcHbK6t1D5TAkgjhOd/RaFGAsrBAJAYccjO+ghHAeOfnCadAIIL9wLB
VL9mlblm7wOUvBJQNd/wW7a4JKwbl9VVZ3BEPC6DXRcTwjGQoBIPScraXNSJtlotEcZxN2j8faRG
Flw7dJEjshs2tPVe9UrS+5DOkjhTUFZ2pZh+d/P8ZgXDiCMaNzTZ1KzTuUYLDbC0FzIkGLvVY7zN
qmKPkuO7DkW00tSRwVctenVZyMww9b9JTM58Z6WMtkLEGqCeANbFfP2rbEnvrqFa/1Re2JHAmTIV
IW1ZI0P//TLc8ZIvUp2xCT+sRyOvX+0rR0XDocbfjjjKVfzPCDLLg6D0jDTb4QXbRpVljUg6jlUn
Xj9S0nGg+2tae8gT4/VPJv1KvOtBapK7fH6z6ED77Wre+2PGVsbZblNbCDiWzs80bw6K8uqSxWyh
+2REzmYi5mN6QQ+L8YFBNvYFrENtGs2NDKpbA3P4bpseaCuqFjdYUQoHnr7dHyCyTrmRxfNUSyXk
TQ7YmNLeMXFx5X8gkCXxa67vJKH9TnU4e0GilADk6QlrArJ0CTUK4LRwI++hQ5w3fgZg7GydC4mq
lldhTVePXsCnrMGQ4YD1USoN7Qh2mP5LkV7o2um3KGbus3g6LuPTNBG9U0KPLP1Hpwr7GglpJJAh
Wc23HNdncapNGUjjqKyPgtzTNOo7ywmR4zbCL98512IeCHKFTyGfOGs3WF0Stw+LXxWGNTSQP60F
ZDdmsAcb16O48uJGcH9EAl03+m11+EoyUx93Jj0MmNRZ/tFJfUlqvE2JducEgS0YtpaUskPFAXor
DLOCrVabOHYjKT2QihQl9wuQtENBdOy9IUCz7weGoWXRfa0nExjNX8WRGZxy7O2dpS3ziz09Z6sf
oLkex6oTuPdhzu6lNDmhmkq9uNZDbVoax6lih/WrLVU3LF5mhQSoQMXDhIEsWX9DdGhrp6DqlaOA
6mw8B5znVfFOowpPdvWU40XSw8cUTZszr0DAgSu1CckE+YnKn06gjbOh8kPYzAOQamEbmMp1imbL
TcNHf9rkbEJ62GvEhSIql3FN2/ATOByeAGelU6/HdyS8+B0b0oUvJfXi+mzw4cGYx4XIO+zf85ih
BoMa3V98ioAyogXYu5K0QjlQEc+rFlv/wKTFrKWuTZpQsb5VA0Orq+4NFBI6wwsJNHIdWbmlMSug
tLX76aXtWlbGUrT1fM0RzMS/aJi4soYukRgBJitkyVp0tbQnTABLD4OLvRPPrI0hYpCxpelAFhwZ
2oUihP9AQ5V61t0P1rB6AoJYqlEZnE84B36Z772TdCK/3rxUiznebO//bxdNco6mioJlcgBDM1uC
XGKsE9SZk1RMAn+stmQk8YQE7r/b95s/WtVuZi++QMqObwWRIUFRP2FIQ4NkHNf6taxrOIvk3Wbd
M39OssOgbrErwmSE8sVS5knAn8Ft5OvxCVafPoEvjim1Y6sP42qBcQyiIH+WUsymn6bKByPTmFfg
AwUhIlQE4I+S9lbCUFH9WLox0DyazqiBBEZVO1mE1BVpdAoAlrrZbJUcTBjU6gdd+gGwiuQSH7N1
rKmvV1lb1Yv6v2sksQLo/JDFkGHYN2DpOkliu7mbpjaOihvCMO5h1/vBqh/BQrw31HnZmhakTslG
GWmb6WB9vGg+FvZn04BDNb5NsNcayGV4dkRLZacvLw5mFQxGw3rcCO+iwJ1pjb1akbNjcuTlNlae
gByQsvlTcgwpU1HGQMPcapwF5Wzv3gWhXlwLnDLYTy7c3AGY8l2dfsOvFPjfO2VaraP9Ktb1Qyu9
G5khXoQL+8H2jJy2w2wiPoZbXf8quin9f1QW8zhrOEU12rUxAlPb7B9BRYVdHBgjy07m7pLoNpN7
CnQttHpk85ftD1+NBXuFMO1WvSK5++sxjELK2EZGu9IxBzgPHVAEks2+g4MB/9bUBPUgBgFyr959
fkTD0F6VNn6cKetXqTf/6ulP2GPKwMhUI6XcRE0eAxsSTUwgXmdkl5WpfLoT5agHptkpYHeuGTco
Jc0aGzbNf0Ar/w9NaXQwWysqp+4yb5Ca9ABA9PVsH9Sd7gseofp+hlRNHswsEydMnHQQZ9XmiWBi
ytJ90rd5N0v31yPboPjZj/Czf598twFWqgRYpGlqjfqKckPjaIsTZdJi04oxkMWaD71UhlPd3rkk
IDh9DeE7Zcq3hk42Qb990K0SBizdkS8+Tz7hxeanSHOvo+ElsuaJoCTz7JlI8NxSzM535NhHsO+K
JtIR0w5plS67mv2v6UPJZevDfomtUzxsZwnSzJHolRdDxmxovmiTXLVr+x4hRP7PMCmsb04xG6wm
g2YD/vmVwBQmir6ZTQHycds8mhR5KqeEgrotE95T00REJlIigEof9xLLS3O3Mqn1h5i1LSmtnHCX
T3mKG3rX2UQUaq1CC3e26I51bGaf7mN0FdLRJiL3XF5El75xWL3AFalvvvRQX/DaSjJhlqUUTQOn
B7gkgLfzggsDykitS9zhJ+shV7TdnBKtji5geFM7lZjU+RGHA5CymSpFxcORvmg71zx0f8rvzwC3
14ADY3dpwQB0Q0GDts/cmhqrxQQBtbtul0eWGQ/+HOjYsazsx04DtV/FW5x0hvN5K5k35cs2FFFo
Vmk8c30s7SwUQpwuexFd0FmDze3qnsfFoSZHZ/stoXs3ZfVyXVBnuFbcXY8lbSF12kkhVmy7CPwS
t3aVUyUbhYUDndWitxXn4f0i8SiF83m5c+xwkt6mIxQUqi21qITEdnw61RhrIerWOX0gCZ1QroPW
F4QMvsAYcGLv599rJk5bcwdiolfZFvyABqavxWzTMtQky7X7Ca49DncQRGh9hfWFWem+HM11V+MY
/IWj4od6b0+bAD6gW9GhJ+So9ZqqUAeiShs75WGHWjK0PoB/e1Xs/1cY4CUPH04MI336su/yiFFf
piNTOD7zdg3iwAlAeYPjKJuviuBJCkda/I21178Imxh8ev++ZOuTUwQJagYThPsgDAeif8lTEWm7
wCF9Ens4AMKmdU/LbInSc772YgF1YM77vwphtrRKxY/LYnBjotyHlK+0kMBTzKpfDLZvuCGAtPCL
INgQ7meTXrynFBXRYdRg1f4Xf4Qb02RR5alyeOB8IM78tvYhmI5Bl8oIOk01JYEkjIWmZvpfvThS
MY0XvOEkuhCKR7cDepHhsf6dR2s9+ZInv8PCtiBcHHW561s+30cxJQ2AWDvQyZTbtjTPXKrbAsXU
GzuFtb2Oen9LAct/fpE1ovCiYxNTdvYS6Ya1USZLuPYXekSPmOX9S6FACkVZyfeDg4MW6mPGReqx
G/Y9LEXQ0IgaiK0r6S5Ct2vxE6EUBs7DCn6kJcHoL/CLZUN2bC5Tc8GXhI2odtfFUJPliYhrPqSz
obscuZGr1a/guWezlL9JFOnJ1wv9/geY3r9F7ELkeZaaMFXWyw0fLwMshS2qS8neF7OHILJQXFlV
+lTngRIUdIdQEBGvLd4TzHIyOeY8lgIAs6ALeAZ4YTMd90MKsDK4ORndPBN58jIx+0g4h55qb+1x
z633HFnkVqpEbXWWRjGumhYqhG7yW1zTZUZiAiHal3lPWZ01NCWFFs1e0KutNZOd6TvNAqZBYIZm
e+1OCYOqOkbnhUIriohMvCRV4R//DwSBPOg/A5cK85F/qzawbbX7bFHi/tsrdNphukio/qPKQr8r
ROSvS09aIPa+YxE4IUJugTDgN+Y1GgD5WYiN46QNPS0bf+ZpeaDpqjgVZIwXgm/exNgFp8K7iApu
vU9IupsXSNCKq0Kfk4WXCN3e5ZsfxGuDrRoLN5o15IQjlLtOd4MaZ3YLWHQ9730A41xWYP5efkhO
9UUsvNbmqYqeeqLeNGks5jOqXU7ug1imvvVv7O47OiVDFGPy0KXnpSQ5RddIrKRtAKFAHBMzspK3
/RtWAzFvjR0U2Sz7Z15Geoi+GHJPTiDoECxmWPPBp1DJSOrxR4nNvEwiqzcI3drNjRgFS38HOaZX
3Sp28psfuC1z0Ijdm5uZBJNN6ez5KHg9ZWREjz/R+tbAqmU9fEyNaviYEnseD2fT6VSLXd+oQ/VA
byiyocjWyjU6c7KgLxNRESKvG/r/L4oiHGlE/n5yRiVLq2M/JgHecqAbBQAX7DXLtMM16W/jz174
B6A5KS8nO1p6EIi4Uy7wUYhzlhKuD7HbnIOPET8MgH79xoix5nwLoV4CTbYZpW432HEzZbXFvHW7
kOKgDpP1UNMD5YhB7zFDS1xhGCigqDuGCDZT1cAObxAroB/ut6an8h72AdQJotnxlr3giL1iChz7
LNWy8CLSGJ+aE/eBMgXyzVAf6aOVLMwnt9MVnT/s53jjUQ2QJ8knFVKtg0c7tIkrNRB3154nhRbP
iuuSJtz8TS2EWJ3Cerybkr6IVeNHsEgom/3V5QDsKedEBCzgWRPxG3bhACJc2ex9PUaWy57Xa4ZX
cUjymVGjf7eq1MdtJohs7M/KoSS/DXKpuVB4+LuISSt9IWOOgkUohpRIHgnhFn5BAKKSurk/jI9k
RvtnOS2oSEP5nGtLSj/24ZMHK2KXmHanSLb10z5UbIUUl7y4ruPhfu6TK37DsXnqTMk5aXOeYGX0
VEL4GXZWqtriyzNAG1fQtSKFa//8XEkP7HXtuObxOIFD6cwosZYL+MNS4EpgmUAUPsCPWoUJfwkt
yGBUpAaU72WEtP5xccdQFMgIKoQ3GE2cBCg2I3jF2/oSydheHHmNp7k03M7E2uHkgfrX+Aa6ctv7
O3PUG3t7sglWBEB2xubYSww7DTddJ3uyfoVs9wTeOE2c5PfrIMlrQfOInDuXY+DNTF1KFLQC9wUp
/MuVW2ygLxSz8G69vyq9QlCbdOLC18eY4tnAWZfrVcisZSOjQFLhohhXNvn+K5UCz9DJtW1fysA6
7zSkRoaEzTLJHhR2CijR/U939x6FT8raGlU8ZqMqBSWNkAsf5wc/grLeRJrKO97ir658nt4wNRy5
swjcU9QGv9IFZSZr10iZxnmQ/ugJqwpBPw0zfsWCzHuw7z0La6aFS8i90MXdCOtNTgCTe71txIM6
qT4tWEeWf1erbji4VPQLRQodkA/aEN6Mi4xceBXonS+1AtjO/Wxt5CiNPGVXNQKIQd2rjj0ekKha
rcVjKCUDcHw8JbYhJEvhjVV/hZ8nM9b1T++B/+sZMIIg7J8yW9rbAcy7n5z/UwgST67UiDQhWCoR
ZsNg7y8qiTlhHnsY+GYra+/r6ei3LnY+QmAP8+i38A7HLTmw27MqjM9fdAgZUpB5agRwldqMNHNA
14woPcGZMb+hhEhLVu1Zh+k4BbNwSTGCrrKIMUrl23hBgCEwk9fxOqeoyyHgdScakSpnKZaKv7TH
FE4ipSGsFV4PW7v8Z1EEvzepoba5u13D9gnoMOCPXRCnxnsE94jTExWTmDgy6xQdygDIlF5dXFVl
N+9iwGvomPLUjHQvE4D6E19hEu73h4lnHyObFT3a1+XAgqV5PvMcKvhVWop5wnQlfoQUZnDFSNYh
3MpMmjUVLs7pip0oNjAEcqRauF3olSGD7f39hkdCB37GxI+nhEs+RbF52a7jae3sT2i90NZTrauP
MI4RGBTrK1ARc/nQ5JgVJfjJj0vfSSLLZ8iGmHSBBkQQc8ZfWWxTK4sLNeOUsmxQoT9KVas/r4PT
BnM+ycoZ0ab9lxt9Bib9S3rITgk2oLk0/iekNHSA/bw4PxWQRtcCAWFJr5npMl+/uKJ38KPHHLja
7zxSNhU19RJ8l7T4cyQm0rjK4uyM7hxP9ns0xnoHVVFS6PeOnyfCY7Nv0eke8zEUS/HJ0IFW4fih
uMF/GvfZPssU5emEo2l7jbjRd3sC/U7/I68mIY0fOmZD5vGmA1lFO5CQcqqzMWvPsqy2rQ6Ll2Tq
/tGWwKkLCQYH9K/iEtUGMD8HiIS9JDZwqMU3kj950qq6AaGcy92vDPJgv3jhFb6F/EETsqrC0cTb
5V79dDsUmY6IaQUsdL/qUAL2xgBXzp/tayb5FMRHB19IVJ9Tdf9HE8he0feJOB7yl6ehAUSy8Nsa
hHf3ed9vkWOvXRoHgfdS983wAI3sgNMVRYqYuX/lTHRmawdvWKMAohCTG9V+qQXFt6GGrQzuvfjL
7556DdToaJdWgjd8AchPUN4A4iQ27tJJm6t1LOBvadYcsv2Owp/9yuueE8YCW8/WNjbFulqR4ZLT
j8m9QRak6JnOus8zjog11P9hFfsyAYKWLKPgmHqpJCEY5AZ2AL8mRLnFVqO+qsJ3sCxjNICwkG34
Hc8dBzySkVyxuCjrmyKH/jK9OiRC2VFiqnZtj7UeSk3K73Bz0/ovL3ab+9SscFFDaaHupy3xSekS
485j6vKdibQD0l9fjFQfluA0IOJCbv53Dp7KiABW068B/LTzUIrpS0l6OmJiWaapiJdMswxs2/v2
22m1u6agEnrqKZufphcUUTjT8DrJCacdjZjF3HyoCPd+fFVT0/sbxLRNoOvgPUdji3gie4JG2SnH
Ruym4cUwoauICrvbCWzuT4zoiibRpZfuqlzec/2weFmpnFugj0p5mMF52FVQZqVWB71b1wdeo/5c
FMkO09iilBypK2ahxO/hFey7guGsQSXPhla8+GaKiEtPirRQ3jviGgJL1Untgp5gRov8899xNq4i
9bJrkLnjQ2m4ksSulG0E8d/BkAlVrnmfuCIhSF6tuWYD30JTUx+vp5w1fyWZzG+600Yz5CDefxOc
oiO27Uv/IsEk2SmC7rSF6RcaD1Hr1RCUDCVqHvWtwvPl81AakIvQonF1mA+LMzYTrjDx+B+s0nYt
OV9Kinne2YKcaQ1ihhlfWM7/3GdMDKYON4lx9UlO0iRDjytMwTzYKf7t0YjSccxTizMdYMTBh1Le
uzLCJwn8exww5Y/u1K1ipedKNXOqW6lxOlhqOXfDEoN/06sDmsNGbV04XRNxGgFqgoZHpoyAQ9tw
Lt9eDYwMM88i6PrdEqKuqDZfth46AgIxAX+iCCiUed5ayjMRrCZ1rWDPpaL4rb/9q1UO/1bKvOle
QnOpINU0KM2i4/v7VpQNlWU1TzOAxe8dTxKdLAewSkiPq5I3bmRPNBv3ClAUQY2SKNeus3hiYGJn
ZzP7P7KqUbf6nQLyL3/Guf3LY1PfzwK3ioikLDfQw74RzV5mx9NgKg747JS1eFSal8wce2CFt1We
GT2KbHL4ozeX94uFl3+GTpmNcT8e9tEwOZdI3YwAkbnBhH5IG89BksudMhjT2xpjgeSVFK4Djg5Y
xUEot+pkE7b23AOG/Rp4tWpJVa1Sh3doYI8R9jqrBE9DoAHxHXcS3IsjZ2TQIVSTQVq7isSFag2I
wUVY3DGPFbAsNAOEvq3N8/Dlov5O5ceiAKgWTSxtJXqr9PXp207GFR5encAaiiSTsAUUsdnINj5S
aU26SNQyc5STxKYI/4UddYo4jgJ10InkToCCnpnJLMSQ3bar8UE0jT1+4Qtv/N1MQBjX35s7Ku3P
zBzq8npctCiomq/KLuQUcNG6rsSlZdysk4lLH8UjfrxKldpDuZ1Tkd6OLygrzWNsyb58WSgYdHiq
IyfBTMLL5S5tL/vrmcqXX19k3E/aO78gohOo8eT+mxFGMike0Fl1sgSgzTgV09wPCBJ31FoOacFS
UeEr7e588MOzkYmQdTCfRCwmkWm7cDZ073U9o6PQfC1ZWmU5CAd2NAxofezbJ9c6uMwhszG1fw0x
/T+y4rpveKFdAm5n7z85e3JOTEPWulkEknnddzl0+XmyyUHol0dsX4zHWPiaFWK403LR/r8LbtTo
rIHBwKTy38pbLvlPSK4hnYbSfa7hHjyxG/F0+7m9J7BCflkcC3IObsdJKWqV282NJtV5x8R3CdfE
kwTnKV9qRWdA16CXG2UMo8gLTnUqcqpu7VqbpdSc6/6zio3y2s3fWjAcEOsJBNLbavGAfSQuguqK
nojuUuhoba/aR34b8R6+LTVdyiGVqtRO4uAqKfoDkgEaIOrnDx3VYBQ+LhQF34YYjVySb0QEgCdT
b9e4C7lF/v4SMfnJpJRJ2mRPeQ0dZbxG5dNxWgM6ebkG/F5kwSZp2ygDazz7JUMhHwb6VCOwxsXc
BaCR2fjx9ZB6EnhOAf6EVxMoi/TYT+eg0wR8mn8mGLM/8xm4vgTwPshOAg2RWFO+2G0hmAhvuOJ5
jznn2ig1/luLkN/TsRJzqDNmaImJGH5cx4XTRaiDIIG4Bbc2AP7UAsNwqDUbwQRK1yyB8WN+USgH
kj0OfH4GbLAEeb2qjR2QQoMRa1piQzH4op9up3vN9tZi0kkYl9n5HYIMUGW1V9KTYEx3wtO1grRQ
w69Tti8uCF2U0EhQCjycEP0R6EVh/zoILVgCKS/y8008Yzqbu3MS88cvvy9XlEz5XN1HT5qMoMDQ
w53erQSypBieKm9unmFqNItE00bIGia6lFaX+Peibnp6QWsyXUzmfNqcQcG9YvvJWPjJw6G/KCKt
yxW6B8eYE7lx4BZ+AT2987OKmC1WWQzCMNu11QkKMRPrefQTZWRmWm6OGQrvk6YEULs9WZcmEM/d
FsOKyuH6iuGH5zaZ8fDGHhgQzbpo1YqIMaph/3v5h7roPxMQUUr0fPZ2C5cjjk9xxmOLULmAH1+L
YxCTJyD5L+dT/bpI07bFfR/BxTvPKGdX6ZYBbYOip43dYXqEKjuqlHUXiQVIY4RaLe2hij2RxH3+
nuFzJOsyGZmHT8VgiSeaJdLtsMUbpLuqsEMVJmzbnI+ZnjJI92LDFsZpV+XeY7OhIiQCkFJJe16Y
7e2S2JTIxTm0SLz0uyYaZoGKjdhxhamebhFX8XAYHm6TxwPDmns+vVdwLXWjHF1Z1JbU+VqgyjPm
jW8EnJFCeJazIkWXWQGPvyW9j5S3CeCCjiqhUifF6x/YBlZmPWjVZjYVnXfuWHIOZP5yR9wAD/9A
/OLRiLegwWNrx+6IC7s+cdzjttLymsP3gxV/6sbkObKrvABnRcykZqd3bC8ybM30r9B1EwILbLcM
2jiZ5d1v3cVkgFA5OGLuUT5lZvflEClkMqLoNAyUfcnDtWWrYgeH4eK0aRALnLAYiGIsr8i11CBQ
MGRQGXbjYzdutrKnXGl6DXpkxqgW8FCjv2X7yDum/2UGPE5/LfwkUl2KvcfHdNzj6YDLuqoVHrkv
LzeBah0Mlpnn6tuAagZX+Fi4llQNjE0eUTtFObpbwixp8lUggqw+rsmFWTb4RQbqTGZT8yvikAaT
SXiJD1TFdmSgPtMG/JMEsE8tj+XZ4gRJ6eNgt/1A2zTT0WN2D46ECfGOf3C9sL9EtHQjdgeQUQZf
MlZcTKMOxrfcxHhPcdFKkoa57SwC6eQZ1uh50nf57jPgr4nbEDMLgezx2tsdkzmdlzT0wz62FbTz
W88Bk0z8aRRvVRNi5suW6ZBCkRtRl9XKZnVJSrqqESrGTeTV11l53k70fiWOshAHmW2gZ4pzNFCN
yx8D47Y7To8DR/R0KVx4jO6a5nFaHzM4yXxj+wpAzOdY9DXn5PqiJKoPyVrSxAC0CoSr5Ekwx2xi
d4Y+wxHD/RhfH2k1C1LxxHZ1Cylftksx/28HRGo2Ja67j9FjlOzl45RSYkWr/vpGrvAjViYvtFYP
dsILY5QqZPghxfsGQL2lG0o+eyTbYSXmCmqi7HZY2ewOxk0SyqBQQLr85zxXEQ8Wa9msBrpAgqas
VYZ7Uy/eZdgV7Q9Tm7PMhOI8hUwbeDKNcyw0AkjmKYv4cMmizkzH6Ijbao71ZVUJmJL36i8Kr2b9
xD7QeDCFQFjxNkG8+Eo1hVShCLaT+fCDuaUlrD+guIizgqHz6kuYRFS98fJuN6NyEpTdWOVe8QKs
Y+sn9+cCihU/HoVor9QFHGJHC5hk0XGmPLWe5oJyrGIviKBGmlokjNXj4bWmansigNEmSVtIzcVn
P1ZdaA9j3v/8J5ieLpew90t1ihFBkHJeDticPqOOb4keWG/9oxX7SZ/jJse4aR819zJmjg3vTanm
FQngRz7IBk9M7EJ+gPUgb7c7oHAAsOPeEPA9tAphzZeo3JPPodfjJHM4zelhvaf9YtSt8O36X9D1
epgIActegXNuJPTvs30PojfTzfZ9m2XU31LfpV+u0/W8zvSEuByR/pDHzXGCHebjw9n+1zHWxHUg
5CBaYwEoZKMKgWtWxqn4YmIqg4TXhISeg3RdFErhGlo68HtOxHscduz4xfHYlGYJan2EYicCfMH2
WyFVfAqzqrkxf9/+oWxGyoJnFc+Umbs/DCrf+P1Eeo5zi82eGhFNXY8mOpJ7/Pdtq3dZ79g2vGoS
Trn6UfhRnd2weiMtQd7sq96uFLxJJ57baftSwilbomBe0K0usmQS/b6mN6Xzt05PLiCbZcI9do+M
EXLpW9TjoMKO18TJcYyLItPdcL4MTq5jINH7w9bNJM+mc+Xkio0Z3EBM1Enz1oTHUKVVF4c9NJuv
7PFQ2iGYFMup+miOB6fh/0B4ETv8PQIz5fS88m0B7/+xXd7ks6QgE9MutUZudhnuTupOzGZ7mE4D
Iq2bbo/gX8UMysn+u0HZHVc24fe8xNkbBfgZw6JTd0KBH8/3iijlROClT88ihxhKnrZjrBKgSz8u
2lNXsQ2iUzZGoM8ll2Ozguha3kW1LlG8dcxgCe+Hbe5rSjuNiMSb/ftoxVrMMxKJX0wZQ57ablL4
pg2Fmoo7Xec9CcbUfc83st2l/ovr85w7si90le3PG1SikHKusAIEUMCoXIMqsRJK/G//p6kTI/6+
il02dHWnauh+zJJfNYfCpeBW8sv69QhemT40TH7kVdT/pJgGZzlpAar5UGe7MSGhAsSfBJIx8z9+
tK4Dy7G0mq23ErxlVY6a2NnOwhIG8o250zIX60EAZr+GReD9yh5ABaZXfEaCLHczL5ijRDQYWvqU
NMJBOGAMnA/p6+Q2gXNS4bGxA0U62IDzbdPJcpo7B2P7Maah/h01xjwnedsJo1i8VZxrRxCgosGE
anVTwkqPX2MeL5uWO79k0t4hgxjYn0rUdMt8NiblpQSIO4MwgHBjJ668LryVlKCM4X416VDsOiCU
mJHh0E8GZ7f1kXWAWM2ndHg2DeazWURJ+OdW/yrmGRQkt340KSuOxvB4cQJR3v5Bm7DuS8/Tjh9e
RFZDS6h7m4VjqUGIMd8S1SyXGsefNuWLCmOm0ify73g1lqXUm9BwjiObICi3ifIRtEuYcNPt+dnz
JYee7aJEIbEHez9HUwYshtPJCMkXVEpqaO94TULisBCitfp6pu1k+esE1CaX0iWORbJfvMF0jF/o
h284cIVz7Za2nweIlIuI7N5Te3bJQiw4K9NK6pC9FPgC7pyP37Jv5tw63/kk2HAhlOL+uC7bTPe3
gRZhZ7zSlLq+IM3iPbLvhAvlz8VAZyb72Qe48FRe/PsHyD+rJYDWqxlodrX554L5r7fBcyuIol/9
h9RjIS/hxLjMGL9ZS6MJCDiBTdSjCwL23LAT51Tnof8BXv2C33QyH94OmDAwPwZNE35Coqg45eYz
b2zmS3ltKqSFTRI76SnnZizkYdci2ZZ7dT8x3fb193yuCJ9a2w2wmGtMLvaql+0Ry6rBv7PCHK8F
0c1366cz33kRyYpyfj+NuJarDWSCz3AT9t1LmhPP+hiLk1U5HYo1N4DYBGJizrJZ+6u2AelduDZX
HQ7ua10R1NS1UmDzX//+soFTLT5daebIErqwoMun9vyzl3kt/wJwO2rFdOE0RyaDQkKO3DE9yESg
f/kRcfFmm0va6ctnXbub121Bfr55BtFuOxFY9cXZ8PnbemsWZGLzHkPV8jA4d7+kPSanSDpbvGRq
rPELajW0Iz1g72EEXwuRBjea+0a4PIJn22dy5htwC8DKQunGiZWC4xO0yHxi3HtFV5wd5W74FGb0
3v2kHWiUcU/vT9L5ngMuiwsWdmhFUI7rE0wkV4dalP1ScSk/46st94hIY/F/2tlQJR3FdQT3BlyL
XjVYfxrPr4uMJ1wmSWrKVslkuY2fztTjrYs+Ig9KicOvjw1kSyDxovpbFCVMK7J7zEcbKjThPyYp
PVsb5iKZGSbiByNC7eaShNMLsrOKFJ126EMCcX4PW5RR7QDvOWKBDA0YOgntpBV/+9gDNUTSb3JF
bNyi9JekNInuQ9PxILtTv/KqJM1SL4UHAy09nPx8EtZ60LvqA6uQ7TVgzFEdM2I1FEwqOm/vARP5
qeK9q9BPNkPKE2mYk6A2K2VZKZqE0t7a3uPqwp/Tz8c93Ota01VdnoEEuXHif/bjFaBWCeWaG6d9
7Tqiw+iy0NmRIb+K8UPRVxvXA0HZZa/AbAUg+1ZaRRceVokpTA6cbBjFVA2lkr135SW6jMby438y
o2ptWIy6JnBoNl5ykeOeU6Z9fjAWEdiAOPIxV/JpFIZ4Aw8oMDwtCfmLtroGWy0n2l7Ol/SAthfP
ROyjLLRK2pbO2VrzfsBxqTo4yUB+386T/CJozEBYCsvZ6bcaDIhLnUhsi33BJ29N4XVwhj8EO3X/
8A8UTRKwRByAcYdJmheB3Eh/xfbHenKPim4uvx2kLHkjmJbi90i/j6uAOL4FYpuaRxGZ1gWGRBcf
rau1HBfLjd4RaSJ/DStfQ4a1a6/1EF76HPmxG5Kt6dbw8FMNrqz24sZK7trjzdmkJXFcwACbdKDz
jpIxElxobzalkOZ3Qg2FnLfpdw+Ex0DyH1rDEODYXImlMa+0SDefsgoVwf180ag1LOFBXU3fysXh
h8OSp3CzKKsYxoYwwm+xxYKunu6vGu4MRsr9uF8m2dRe2Q7ZISX+lEOSejeDZY3/mJUXMYMs+rCk
irpTYCe4ArUKeY+ueVi9R73rRRftLLpaXlAYwfgDQ16w8eaS1F3dmOS+OgkLwUIo8CwT7yT8Pe2s
fS7MlPNTUQ0/Xg0yDHb7/7NL10JI79ZCdjxTYQEMa0DQpSij8jdchwOuFPIq56XBGdJpQqKQCOhh
8TnWMszuiD8UAQOVBTLX98sSvNKtlG9WdbukHHnVYHqaUZzY7vbNwz6RuNHi1gKwVw4hBwcgI3Bv
YHfl5UGmyCSUD/SCik+QpUh39QYfJ5mra0sVpbDDsx82k0xeHsosr+Le0FhQ9dgYWtw6YFFP6cWa
ViCpVmd86PaBv4wMSPmR7h8cBjIZNhCAgIuNoKPnrVVGgAInDOLnpjk0MZz02E3dcHQfcdDHSCtX
nii1Ncxmz+Bmbr8sTcAayZB3x9Y9MAUbfp0yzDla/FVXj3YOCvkiNsThuSzeMikhS95grpY1c5OH
5EKdbcxHNY2n8fGUWSsrJ/NvBOEm6yDj1CTbXssJd/z436Rvcs1jKCVWrKW8pDiCfSKBnVzO3hsv
IDSp+StFWKlpChB/nrtp8R4wslZWnfsTWcW5F/JJ8eW7N4gy5T0H5glQdK3S6n8zz8rZgEC+KFjr
1uT5JLYrYUgOnDlIPGZcYt/Ri1KmkDHTAEyXdXeyvM1wL9p/2AkGh153PL1DOCcQMY4GBwNy9Z7/
kNgjfPl8jnzpoDQtIGcm0hF6wsSqFi52ytfBH+BTwZdvQyJcXvUKNgvMHBIbaklrd+HngLrNXZOe
ttPNkOUblsIKaZsUeevW2JOF8k/FFQMEhjlsFtd3qVEh7/Eu2Vn0p8QGr0oi5TV0imcWr36cPhYV
vr82WYrE+Scs8yWiB3vwoD+bk1zCysZdy9AfjNHWsZgh5ixqaJ9xvbbtXNvvp+NVdiIYgY6HEUPc
ipr2SAp+yeMejwPKI3U2E4k9Uj2BwSMF0N9yfkV4MEl/GCwJ3maoC/KPBuIE59K1umE3LVvy7Jb0
43WvPtbu7EQiUP8joGif9JdGUylrXNYfudetUo4OE2fcJsN5RwJOegC0fD8mOQ+DHt77FzNh10xm
n5pmTvsqUmw8XaHt5nde4mzPZyf87hXMA3c1obrgQf4lqWBPLYr+aPTBq3D1BWesOi1SMqOlDHJt
bFFrklqBaXZCWRq6ZG3rk6g9ItZW66ZwEO5DHb2rX7vfwQKECjfgvH+cvqTtQgbyp+EXzt3xGuWd
SjaRZqW/U4hKbMRfHClRZPxyMUJn6bjfgmuzGn6B2f9E+HUzF4eKzJ+b3uXxsz3/cg65sYUkWBf5
zvqpcmFwEtpOpqfeB03xvsOugiJ/NfIm2rEZmJE+JWMkh+ORDVDXYs+WckhyRv8Bi+ppHAvhPDZU
0EijiJgsz9ADpmgKH3b5mjIr+9Rgz9I8h+Q533XANN1zcRN9J4NqpfK8Qg8EoO5U3LPjzfN36YLg
oSYnZIzMyena/5lbgNLDB+vUAQF4Cuej7uwcWztmR+HX9W74H2xGlKkV4vEcjdV6WWk71B2o0LPU
OT7hADFh+MLY8iH4X5nPEAlX8EO91quuqbxg88DRz/F0sYRP/weedfyFo7J9ZJ/fgeCWwDP1HGnJ
2vYNY0+c3dUTQNoEOAV9no2cCZDllAVq7Wcy20Ez/QCCxUsLnQTwri9E4Cohs8cdDtXhHtxnnIKN
LRsRxXKrv0E+phmaE+F1p+CoceCPQfp105dH2dnTR6uif8ZwA2zaK0VFK2vjYHlS+SVDR4bIZT3v
xTe/bBWaT3vFhgWolV9Ki3O5gX1b+N8Tzlv2TuaKDwrRzlMNXi6PN7WfC2/rZSYsJkN58k+/9r6O
/nRJJkrelRLnnsmh/XAy8nL+IbOr7EPJYEW/kZIkLEHXszKqarCkBBmfOS87+QXF/0lHqkOpfUSb
lhoo8Nc0NmEM3IKZMdvP1mN21DJbrHYk0RbAJGHT8yQVzHT4BjKJfC0eUKi47xHJ9oIw+TNhLEPg
G3pFQlP/84jKel6sxNIsN2f/z8AK/qwp+uiIA4JXfFOKLsCk3X3JryFiikBlC3HKTxX6UaQwHBt/
LOqqORbxcNQd+bU24hf31gBj0toJkaFn1I5cf8JeFMN5tApY1+/l2HcV1zBvm6MsvPo1WuozyqJ2
ZTxVspttT/xj9ZzXIovFnxIMdA5gRUYXgjM7yJkwKHoB54K4iVZezllauPUiWeR3POZBBJlE0cue
msI7hkq8HwVnAHY/90g7wfcKKkcKaN18EbExDUSfTCZqOfzT6QvPWzuk/EEEmLDWh11sxVbg4JFB
cF3YMmLgrciMok7bS3lniemy5XDPhe/BYx842Q3WVRlpffGk5mX1xEjNxf4a+0869fzGAkdQintN
RfsJw1YZ9X/lfwys8vGHgUmcQKNeRc1CWIOFL4AAYCG3NWFIUFD5AYAYCjFHpg89CNu5QKgMeVr6
LayqG08aWRy3cNW98mfbOUWMCcg2G/qZr+iAZIWLhTo8d7aA03SUjbFKakYW9p0pbRm5dvkBLkQA
5zyyegGCT4rcMmr3vT4/sCdazW34/afKKoLuNe16+sP7n1FSZpfkhLS33DiXkap2FPTbHQYDKZt/
8mZUJDnm9jUjqskIRgrbHIzMqCXxPZJpWnRX64hgh1iRKwBOuPghrojqf9EIzESAZCSmqBcuWSUi
bENpZQyUUth5KtEdgLq0LUScu3GuX7ahZXY8VhTywTo81S+Oa54iFe66mmxIi/a51tR+fR56rDkL
mRh2LLAPgaJFtFdmzyJQZzgfLLUvHyh1lkgUK6V0XjOcNpGlA4hFz1HQFuk7/PpbKZ/28qIb7bhz
H0VZduuLQPREMFl4+kOxl3olCOGFZprcJJmbFCz5XLWvjF3hAGMpGmpn680ah3MvBgDkt/VoxXfh
YC1QXW4IriXDs0DGc63M/c8TMqRpHsk+MDP+gcL+gkQH7QPn0YDMDVHwVYYsYzTMYDyTGJ0a9T3A
L8uVhlyhFJYIgSEvciFBzRusNFRC7xes991vViPed0t7P9ZVRJzKF8SJ9nL/yYzlXFU8LcxT1iIv
vs+ESdH+/rSalUWlB2lOAfptM6jZyhc5oWhgMH6msKs7WsonKlfkN7c4AiKY1tTrjo8Xa6AG35m7
h6nK16tmF1vf2euJZmCal/8fYcWL/uDW2+kPeHp+n/Yh/3CAzetn0Fx8xWomDNhxnspgaeEsb3Kq
kzwQx1uL4oLD6twvpFtRh45Fvahd8J25qj4z35+uC3zozFqhHGlsJEoU2MJPGqvsVm7GKONyVs2v
MiKiC5DZb5t3p17yUNRjAdMYy9iCNWsOd0SAfgVzWS83AmXj1XQwRp5u5OYR2f7xOQtL/+8z/88x
4+kg59w8mZ76i4z6N0ZZecpbJdXBeWRcsy2y8McALIqf0N/dpYmFtAmfPMWA6+WunAl8CDeQSTZh
1gyJc6AiMsxxvNl+XvSlf9Bg61AZxcVqdDRDalHRu8x1iIt0TC1QWcNfPLlXOkPUTXV3Llu6qKSA
pOPN/xOSiq1HgwgnIZ1gfCq7ZsMTN9ff3Ba687c52txKsBUMiHPNSmYlk3mkyU2Ob6EmUScCOZpp
tO1lbFUSuX2sel1oYrl6GC+oQ4gnsbKNd+E9ImBUt1JQBT8X0qaF3T4/0cMhrwNWIKWpmbcz6aug
dJIQdqf2U73WZwrE87Y/cqhW/n1mobbwnEbEtOcC5TFilwneTHPGx+gbIgsOIwcSkZMaM3L9Q0W8
OMJreLR5uugcXjF1caTtQ2SPq5hM2Fk7KH4FUvPLeSNr0Qxxth3Nbcvjxos6Dr08/ldV3nZxzAju
XMMC1VcQQKMAGCW2GSLMkoPQRFuOuFC6nYEESCFEVOq2jdO8EPgWZq9B84MQVwfm8uCfHSdv+mbD
QRJ0TJryXmnGmDu7PAS7O7WY5fx/EUZYwYzWs6PFtAuqygOruwhWBBShY7r/uarAS/Qmclp10LZf
EyfMrie3b9cKR6Qp0DQ9PZVgx9sMKZ0lacw6Ba+FrHkeCgOYnFmO2bBBYC8o1xqFMw9V5mNC5V9K
msoE0OjWWM8PStuNet62mlJ+UTHmTCsZN678BUGVExYFlRAQ/xONAK6ZP+L2H8aSUlWsgBMACE9J
4D7HBVrD0tdIIloj4NUe0R7lvkhdfWITmbDY/esZ4cSGu34tlyFUaf9IwVeaF39jZ89mrp2YV/kC
tbBjD+h3cCtLQfI7q18nAAVWcRlp+cXXkdKbwOo8S2AhWTpQU8x5t1NJsC51whqxabw7q2u00e8k
zW1LHF9/7UueZo9YYqjXsOSmpFTPjbfN3gwFXlpGDNMV1h/c0Ht86vwAAdqwYYqQFAQtn+K49GMe
fyQnQ5jtfbd6sW+WcBudiFIIa9u31vGoNC5xXz03y33KKws2JqXTvoSS+roKT/uJLn8y83G9gn/L
7rZreaxBfw7dQnfRcETSvcDIk9E+7NElXCCGHxVFwaqmS0CKY4LjvJlcqpEFShA9JmX2ZK/anyqt
xENwBPUvnvI0vyB7LnzojkHiuTUdx5EeL104lUKsayWehCW7pIkUgZCqSX4zTPmOxAU3Oj0mkl5Y
pH7pnWxm3E5/nx16/swiyxbYM8vIyA+tNbmXFa+QleNdYQxlddutnGb0wJn8Ii9hgQglogBdpHPZ
i+G/xFUBCkmgvRQIPGViBqw4ONyaycyakgLjGU6WqwChc9Hh+gyQoLrt74UKspG8gZ3CMTouz2fP
xYuFK+oiVVEfTB5qxJmxUF2L7PiID+i0gUUCrUa1/I7utvddg4SQshkUhgp8Q7Hnkg6j7tNTwBfQ
q/940OwBbegcjMl32PtG+rNMf3seZl+L8y9Wk5ExzPSd0ttQlEXyLcI1IAsFQCl8z1WwMfVCJm9k
aF0L129Hlz/a+5Fs2QvMB+Z+UgLcHZHHarrxaDmTi3x2OhEFITwlnKAnAmVuGUvWp3rWutGuHWcG
HZCpuXvUuyvnnal0LqAEy7Ln9Czo3dN3JiWP4m7CRZdvhWrmfTIcVNBkRypqjOakMdaQC9MayrtU
mYSVSFM50u5ggDM96r2zsejsN5r2jTk6rpC18GXX4cDWPpW8xTMEqMO5aYj/L9U9a2Diw+HeujoS
bxCr5MAs5XJ4BkEggfVZp59kypV3oF4ft6HkVt6IF7RklVKhX70zKuBx2UIieuI4SUeHn7hgIJxk
Ay3frIg8yYL3S5ROcZ7l4DIF25NYXRMmxgyRTGmwjqdVprfSb2cNYKhUkeRsBuvoWSEii1ZY1UX8
+XGeerO98hmkWu0oJFHueNpDpdYz4vXcCbiKrio/aeU+pRwyEDblfPoPu0CPqll24oSC/qiTutZ7
isxlOzvDKDCJAEKoAjW+UqdHVR22ciSd0Pm7w0REGygspNFFYDdzS2N/44Z9hTTbl7eT2NsH+PJJ
P+Xa1S4Y8rt6PnNSQSFHMZfDS8+ZxXkRWgTgqA8mxsQDNBcYRm3RKOPq9glFGEwBlNvgiFJIZL0d
W7X4vwFWkEI2GKnjbQImBFudvzJaHmGBGizeFkUE2plRcO2qSjE3bz065zl/Y/Dyse6PmMB2mn7z
d7kmRZPXjdOa2cifXLaQeCF+o6xv4wFOI68sGfVzTZxED5ESCah8rf4HOX9kQyCDO9Q2MMSn2C5B
zj4t7EUDv4OHa3jXa5FFnMgsX2lq21qWzZKBA2I0/8XOHa+9Gxaxb3Dtg2iTk0qCxpsizjXNjHsj
aPSk4UGVSU/pFGUb8DG/MT1+Im2LNvDvlEUv9VhdlXgDTabCzF0erENeEsmjBYUAoHF4iTj88Eu6
KhhQxf+dXJIEBFGkXC1ZzgTDVexs4TnYoleFFmXXbPwC+bYfsLLFKyco7jHFk8h7/diJ8gAEFhi+
6hEjD7r7GAHxKrI9iNvEIpg6ozG/s5a5GNNCwUdF/RB61wgpIXcy51hAmpH7UEA2RDxrJGlVHrI4
+AkcO5PAO6X6dkZcFVldKIXaoOvvsfiXLBBlRdgDqsGMnbRsPJ68wsUVL6pH/cNq+m1RE0xILaf2
zd+lkVfeId2gaxidPZzZWqotpDwowOgXT5Ja3XwLS/3q7BypWzCxvToTuOD5Y03ZPfNtIRSJ6WEy
BxeWBdoE+juzZAPG7tTJCauCsz79gXmPG2PC62scQ20g3olqvSgRpQ5CwaxY9YE/eLq0tGhUXtDY
DJ4K0QfsgdgdGkZY8oF8ntM9iIbrPaNgxJMsUkdNHMag9+1tuTDc1Ojy+w3r/Dw3Q91/NKwF5qGF
yyoB2751cs+jk47ox/+ySVKLw9gCQ1iBMGr9WUronBqQC/3dNTHGAJ36v7kqsPBLcaqwwQT+X5Sy
SljScNOM7/flYTNqxmeRBSUHIdQQYgNq6hbBY857w/drIqq6P/HUQPLW/VRAkVMFKbySaCTpnaTO
p5TKd5KjHU87BN9m91IXv7HK3PLNTayADzK44kjhg05IyGpEPwp7NebcmVHE+fjVjbBM9SWQADJk
JScdqa6246L8CgMSRiPP0TovSXZz0nJqa2ISnTOzHtTqp2DXoOreSit7GYR66hRGfC4O2slfUGv5
nibdNoLYMHWPYojOD/sGa+jujxY93tSTyX7Egu5TiZ1b5GSCr0IaTeMWYgWa6TxNoxfTMrnJHm8r
uqQ2qqr1nx7jsD6HXltzUaUFlAGubA9pwZ7QC1PfPklbck4FeTEhfYwR68Pb+cd8U7QDVTLM+tgC
cWJQck4vRmrbGM+bAlPTuOTDX1FKNmY5647H/QtPktb9ODtdWWU15a0ybYgAuoyKEUNO9TzBGBOg
a7V/V9sjM91+dA+iAySx4+4HxbehCMH4/jt9spO3daZqXoKD1js+d9Mf26ojzRrkAzHqunOg1roG
BSq9+fmDmTq7e6rIIp6G8Sa90x9Id/mr82YMv21uxRaFp1P9nMzZQcO1M7wmG6319SkdqLQYOblM
sZaPkOGRCIPEcb4CDc6VYZO43b7IOj0mq/IBxfA10R06hfjPW5fRmJlR4iWCUx9yVKzhoFd07YAh
odKzqz7ljws7ZfA05n+DEzZ23XN7sqCNmERE9qoHxc2a018Zncv9PQBZnfGNWuNSqmp6fi9T6NcE
HJabmbSZqI9M2J/efxjFaQ5+7ZBa1gvNR4KPeWZPNTWumDDp4mARYm86cYQkmBFgDfNlfjci3Y3A
es2gEoW0OXV5ZfVLIz2iH31ZCnmQmBU/QA5ztSSUtiafcKdqi/S/04xLfhhwO75hUJMa+O6gWQZX
MClstCCp01YJ2tEhupo3DuWAIiKMjMSFm4OyDUrm+fm8oyZwdLn8DFhMuDktPEr4qKHgyRTx/w9R
vEGzEkuhxYKwkxe1fiteVnQRaX4jNs38dqEWNAYJjV/KgqxppseHpDsYojWODkMsyTcZv9fcZbqM
KizuCzJWTCD0DiEGy3XtrTgKF48ODrmGbXcl5MtfVJZFHqbggUiVLzW1apwuR8wlJRFXJXEdf3AO
cRh2ep8REa+3XTP/ysYijX3QCZKblpdMeJIvt4KXqqBUMwb2RPuciV5hph48toWB4SgTf5FIJ4HH
MdaJRAQi7DYzyVzgGFspedQWAXE49OaBHdY1fX6trqyLm/PIm6nIAxhvQq2Wwg7PF6yev/MC9k+j
COtW7h/bWi4APjhVXsXT0Ewf3bFDQ1HTO9/rLiCvwYEq0JOl0Oeay3dTvct+uC4De3bRc1jGax6P
RzNIPanJa6bGYQheBCkon8HdxgvEm8Qs1/GU8QXgMU1yF/bUwDVTpq5VsmXF/WUJwhewIUYQ3yi5
ZcxPrue36mCM/VDl35XJY1hQqEaBv4GlgdZT4r4N+Wz7u/7o6px8esX+xPaOplbX7HqR6v2/uuQy
xD/xzWQRqbxJUwdawUvjr/mXNrfzn8XEb/VQ5w9cC9l/eGVB8Y6oAr+VfsAgFemZrrBWkmMYLwDE
wwxV7U/1hKzT/wNLPD2/p4AOcWIsmZd6JgXobnPvLN6Xopx/6jhXvTH4UiaX0Qbdyi2FgG2xH6FG
C2v79FOl+XcXCzsXufoaslexsMIjs2jVVVhiRP7pGSkOsoorRfTezcQVDJd+SL8nzKhfrmo0epiF
y9wfSmnjMKDrtR+V0f6OOMUhOs8EWuspgcH3jEVeECr4oezgOhuaoIKsJWwp4ZG0SUBZmkNhMQ+C
4I0vyIN2z5UpwQgFlaLOgeIm+bPawj6QxDWrFmCFx7zsRJmdANYAiYGyslTSYzTySzCCwL47QqFr
2786NJElY5NuKHg1kix87QgE9AVGzMxOUSE+ikJLZre/bc4zi4K7svAqPw6dkg28EPoPcl3MnmOf
Y4D6eks2s0IbG6y1X7otzdCEa5gbEzcaqkJpxyTuzYeijE4CGKYflczZOJnEl03j31eA5RAHC294
av0IaT4ouJNHRsmRmh/kUxvu6nqsPKccsxjao/8WqAya7FvKj8uATuFOGB9FM8wt1yu/fofYAax+
noxJaPZqsClx0EcUjN7RV1RI0gQ257BoTrVqXSTt/Mm1PR4CMnLKd/oncF7rwsSz9ALYGEajloRd
Ik2ZWzpwMz8E4Ue2lKAs07F7NC2OO19IQmaygbBlWBaeNPHi+nWegvoTn6+rPXSXvhHQtIZBBZyi
fTQCo+GrUH1Ly8W9a9Ytk/IquiCKyTb9FV6kj1Iq1hCIokPrba2vYFUWNfiqgU0RJrMuXlujFmet
gunPdZU7dmOK7JkPezD80YnV0X5ZbDHQB2mmPYmfNvpSpyrg3W6x33Tz3lb3FWk4o+ugIY8zSqH2
W0H37yIHP5VCL9StwES7k52SYn6YoKdY1x9tISKpGsC078ghgsDairby4PI6lwDBHBTc72Fse93T
SkimscsZlBeP41GBkI5AAxh+EM+6AHtTLBjl85RWuku8fWV5DoSMObvY659tVGGVus3T/FlN+9bm
huJnUpqiRlIbQcgqryZbVkdqZlD1qFSQikQFCX6jViwO9oJ3v1B6SshOQMOWEEvkjqli5q0tTUlC
LQsNsgI6RyWUU4hsvLyuR43bnLvvyVQqoqaA0OON2WYW/Vdcq0xFYdxZhpVSlc09C/t+zL7bxCio
jJ9YXSW31i0T2vV1GwokDNaiFKnB1RyVpW9HFTFmAwRf/rMCCyV2iTX1+LkUiH52osy4LCm9lmhr
/iIhys+GRFJWOPzGZIQnZODvsht3Dp5qIJem8DPNmNsJteNFPnae+LmobH0YLPyk9w3Ycoy+1XGX
vLYFx5wn/emQMZwYYoVZMOQ0Q6XdchFmq8F0Fp1PpPadCczJ+ompvM7Qpow3+HjTj73tksCN77kF
iF/kxY0Rs7/2RewRiYV9EduEd9+L7/z27QOO7KLfv3OCfPDwKp6fx+b1O0ugvAKffwJ9IuQFahO1
1gU/03wePP/cnwt6gclSPeNJ0CM+z8xMSJawL2+ttVXconkLtdXmo4LeD3jhYRk/v9VE5i551PO+
3t03il0bOlo5ebOKA8htIxTyuc6JNoQ2e1DGPs5O1lV+odzsf6xOdw9x2xpfJQ9kj17avzISC/LE
BTmzxb1+e0uk/stvsUAwwXLMP6hNgASb/XbDT2H5u+m2GJIPYrE1AjUnvrxEvMwtcCtIDWgYdqv8
uzKTdp9Hdwi8de5TAxv120O4gH1uLUdsHoVqjX0RmnK0uChXmHmaIMlNxum1P43Pi0iKzTtGOtsU
Cz5LXUEflyoV5uEz1hprclsBnnhArhSUOLciLSzxtfY6eS6WWI0buxINRWm+PqjpClXDrteKeJbM
A5LhBvAYXm4hwVVCBBZd+PAov3XzSVUX4w0brWC6b/sS+z9hk21d7JlIOK+WtiZz9a8OeDFtKR52
YbavM3uzG9hmK5LkOBZ1e6mA3qQE7hF8dXZM0OcY/Uzx8c44QHOKYdJty+77gvieAQjd35kbpUoq
ZaJ31d8vaKXdjByTDPWkXGq74xUkMdh4yxWIcP46TUZ4ViRL51Fg/BE7ItnuKXMrd+g5ck3+1BQq
WzSQQXfpZm2dXdflaiuqRBHuXQi4F2hcWoREoDJU5+kbfvla/dLXSHn2yBh5qiXsUx/reIAmaCzE
YfipR8tTOFQ7H7ZiC6wDg7zmocaBoQ0IbqpLB+3fA8XOAtjzqcIHQgpMW0K0eyG43GANkUB3EMkZ
1tfdQzghVbyXePUYHMbsCqUPvSi9IGRrR2o514TYEynTZN16vTbLwg9CK5Dh46SphIXHYwOgS3HN
y3akhDYIs+7STnZpiT9H9qhuA0WWXz9KniZNWQXiA56rj/QNLv0yimJ70keFt1rZSHyMtqHMRL9B
Hbm0e37XK89PB9AeUVMKckwgAsAQ/PecyFWCSMB3bUES6dPCdXagXNtNaiUsiPov2UxGDhs4HNd3
XqO9zjuQY+rUxYhea3q27bbzZA4AwkoPUtUE4Un1ivg4mZ+OqQ6qi70qTyihVWyxjywZVMNQk6jR
zL3Ifm6yLEoKw3gNwsThL35ApIcekMUGjkRJY1NSFfaAYpbhAEoSbIIvYJTHeA7UR2omuEt2Mb+M
xOoh6ocmlWqAm7pi9A+au4vjGG/ZCDvQf+zcWgctu16fuCp5Tfix+9p1g5S75SDUVmQh0ssF43CX
3qA4/lbnCoWHEHrPpfs0j91e4gy3qBddcMUV4/RFEqcmT0n+JaPHlDhIim151cH/NhbzjfTAZFbO
ClrmjwGAyTOkKxea/VqO22u/a31xLkz77HVmmtaIn3kjKYc6WAc2ymrC7W3vVyF+tWIwOXvbXV6f
OUIHfPPhdA6NYsya7SzvLc/YNdE1T6CZVEayJaLJ28uGMxUSCwqff7RHXAKLePNm20hEn+Ir1ik5
5leoAjtwn5J04AHTR/2c3I/J1Doh3UT7bZipyoqUgFuurg0vfSU8cN9gvXjqkJQ5HccMGpTp+/cP
ND5wvraiRs/2TFRol1RSJE7IauHJUD+QGSyfQGRBKkuJZ7XOCxRDyVhOccHv8KIdOAGy7F78VxB9
33XP+BNUJcoVFabza4CDAAmaWaO1QB66iPxdaGlpqKQwycmBlH/4QcLfgQ6zDz3icklUDT44jSuz
oZfGxba6IMlltO1u9550+976LE3fu8XIKbzXNcAsqHmeEctQ1rgIielQrDL/AAn6wnWpWILGqChp
pZG16HKIPS8JEedbJpnPIISowtlIbUu07mfRn89bgCEJ3MI8BwVclH02WhIFxj9DJS6ENwG8fCfg
BRG0WM6qAnPgpqOpbwA1NHkH+lIKBHYN4hZS2Ibh32YNJW+elFOvZpwwWPgS6farx5d82NDkQHS6
5IZxgg4asA+lVVme4KjzsZ/1Rpwd/FupZ2QAO+LLZ479ryu+fMqaH6RlXc9jX7yumCDqEO1t/UfF
7all6pe6jEOlJiC132vaYuT1j1eJVTcIZcTtF6YkvMTm8jKLT3CgAJh0YW49WkOq2qAXR5oG9gQe
2VuVwQkiEys5gXY/836F/LiB+w5jN923NUU3udDginS1FHMe1yqPYNy+O7XUiFpsgOUMDMFPlwFO
FpozcSVPZ84I3qA3WxnNU4Jcj6DuTerIo2+UFy4ieUjAwtnQF8zc+6NOBFvRMwBLs+i10XH+jlq3
BSfwWSaE0raPsnQlxhooN14C1QNiO22nCTAsOd5O0OYEF7+yHCHRGyFN8YNSrsCwebjuC0WnwywI
3y2gLEh1mjdOnHFDrTQtA5I4hTkNaZWRTZedgLB57CRfi6m5MrtsB8cWCQe10/4iELBWD/j/2Us/
SRYvBZfYw+2SBDXrYo1ZGjRrc0C5dP/jy0fFjTIVtv5aTt1BNAez4Ow8RnVXDThO8XSb0BTzgEMs
9do9fhsknlXZPGH4rzH1Wb+4iHP2IUePH4FBOl/AIlxLEUH03f2n5BlAbbe/3Da3wM86hTSvHWK8
ctyQ7lnYrSDM49O9imqvlF5hSq9Lu7v8A6H3kAeoqjz2angbC8B5Mtyon2OOOx8L746gdi+fTXLC
XErMlQDbKYuVBKj977bFLecYIJMwdNsQ4eyrnWYxnBoMl5z8++i5+KIL6z5kv6ydAog2Tgo8x7fE
UAPzRNTFuMrX0sjbxGtzHlSg+ZXBGvga+xGToXwjYDkLRzDMvhBnKljen6EYktUn+aPo53mXnHcR
7krskUwnpNy/P3QYE/Nz8xXWfyUd7BTNQafA+s55FljVz6LJ4STyLCz2zCjpqFMiZDt8P5ryXLHt
dMHyCG977fgJVYZ3MD/SxZpmvBMiUw7RVwvr2FrrXD3q34Yv1XhbDzIcZkkhyGALqtHD/MUaNFGf
N45UgXSO/S2A2ilsoFN8R6wwJW4osRtgrwfNLarnT52wj7pYbTH4fubPhpSm0w6cz5vvu4oZJ8io
8PzPBXZ3SVhz/B2uSo0yL67ych4iUMyMv9nqaqUN1POd4qlQb6YBMzISuzuU2xkUjLnPav524Ec9
Ovh98+EYKzzYSW4ytE1/bMmTfR+Tf8/hOy5BLZH0DK+U3N7ik7vpxdFmNON10xMTRRHydyE8IH1N
4mjgK80/fRoknkpg9o4VOI2GryNXWhUFna7KvAjEcl4yiZL8J/QS8gHCfHKCZjJyHLJGXPmJv69S
A7kPQcCBxJJBGED90bJJ3Rr5hXi1i4Q9tAbos+LVmaGVch8mgppY7vzTvJZxiagofSp0eHd3779v
qTb7qQyAUKJVSR3GoZQe2APQ+t1sA9k6LbTdiR1Ni5HxQfm2o6cXHDUWMLRJvZSK6STrIERu4sEj
P27PAJ4/IxTeLv1TD4Gw2R9Fl74/E1i4xjrZ/znlmZjeiX4tmbaB5eyNOcAP8RBhLoBemBwocpZb
IppThwLjo9YHyOqEda71TnkCRT+765QVKifq8qiCT+3qT9WOHMsPKKLHV+5jq5O8dPTck9omk1t/
lBxYulSh/0WRHxbMi20DpiUUuhz4dbjUe2c4G0OWmGwOCsFhBnRbtiThvFzEl/fgRqhJONDsRQga
SVvbc03ykdFZLt0nydWZSGqPrw3gTls7nPjZ6J2FTGrXopZo/8PTGbimvy889PhXp+e52T8dI6lP
Z+JWTBCRFClLFwrg/xeRUVBRGCr1Uch4fIcn+V5m2XZ+yVqL3OK5n/6Vva9kGguWAxelATbLYvYy
3q5EvyvU9M/LkCFahI5YSuS/jTEB3GfCltl2smDYZDRf/hmgjhc516lJdHmGxd9duRm27oO6lxDe
yapm0fSlAdERrk+FQK4RYy0arTbA3xi1jPvAX7JtkadAZ6YGSIQ2n4siHtr1vDnaYWAN/j2lx7bz
0Smtp1h+BGD9WAvQEKrU+73IJua15Kb9U25caMGZnKoE4n2Q8wB/Xix4HdssGb8qfuzNJru1v15L
L7FEdt/kZxTPGPO5QL5/VyhtBazhRg7wyvjlalxnb55pByc6h4TUm7TqItXk2tDIjiAoQyYMYZ3F
AeJ0josWR2WimRDYycM17MFkscIBhoYRvtDEMnBU/FEblMitCkHasVj6SCdQpXBtmlDHE1jTLaf8
vy+gQGDp+yDtT/rN9UgjjnR81vRtHKwx14fEH6zPb8NjM9142FiiZhvg8P2D7wBTv6cxMGp4mx94
NhlgU0rXA0UHnDBZFdUv6hXihWhwrj9UOCm0XQxtF8UCUdU6StoJ0/GzTleiJXQTFXXVpdTfR02q
admENozi3PvzYv1YeFRsoh6ssJ9xH85fCe7oSSB/w8rTODbo0lNYSuAREUkqcIlrXsE8h5MEWvIz
/sYoSBC3WW+MATv125Jrduu8FZe2dlvmVWxuHGgnkxDFoXjLJwRk4YkYMhRy++Tl0qyThFSKntbF
3z5F7YJ2uCeB0KINa2oylt077b+WRPlYz875stDMBOT/xg9oGvYnLxlEv3GDitYRf2e0oJiJeUUA
8rz95cSi6YFi+FYlXSCDaK2n8P1/ud71SFeqOjnfOC9h+oyB4dHtopqD4rb9NogBpqRUFvbzhOc0
YZUvEqTDRxsIDe8ZYbifqWv4iBw8Pxvmx4FrwSGfQzEO8c2rJgimGV2NnKorKUYlz7FgpykHJ9zk
W10WgH9C7rdcoiJX4HZlwyUp45YoC8JgQAd7GQgOHj4f8rkKlQgMN4zeDn+Ho9GMyS1KC8RpWFfK
K/miPnk3RUqcBPzJofwbWtfrKEYtlTybAiLuDn61XUZVn1bjM6y1igQyVrppYKpqhiApzQyXxdGB
49CpimO+AKDpCLJ8nJuQkeO6od084Ufj/ExAhtpBDK7ZO09AjvwnO88P7MgDGzzA6Ps74Fs8WysX
ThC0TfK5TsCVnIHAgO0Ug+LC5W1iV3+EaR7ekb66bEfbp9DmD5FeHVFFcMvgp8k7ZOv/4aX759Ep
PWw8b6LUCeMhJT1HDaEY0Tk397cuVRaHAGGzGtI1CXmkbu4xoLT3hJ0xGpmPCwxGlZ6gCdLtyeGa
TtL7ucMrHqq0Ejx42MMgH4JrD1FnLK/J3j/xX+IA+sSZeRyUQS/ocZaQHWwwUE2epm9oMZtNxdTi
B6cUpm+YodTfaIC8V2UDJ4T3ukZR2nxh9pwu+d+5IGMWZrEmQFh5lLVczHvRiHZVZ2wF+w2FdHmC
GDPep/uYTbUUwV5aF8bSzzsCsRTD0IV/8LqUOAV5GlGw6yBMjq54AJDanIq76uyKLlm8eDhZ7cVT
rkHmr5g1vpcxhTxnnqDJLfdyzDLwVI+qSC/FXyoVVAn7/UUOw4/uOnVJfXVunQMlIksz7hzNbv7p
33SKpA7KI94QsXKi5brfwy8QrlUIbabVbi4FYbshBA7PuWas9h1htSFnGgG+gwgXtviKRKRAnND1
hp5EHbHbbsol3ZJ92COu59uo+8HxscE2AisxnmPce8A/Q6x0wxw/R9MSRABPqcMqAxVa5Pde6ZKZ
3fQ13ZlDCzBJxR+e5I96hBBZsRgSZriBmkSnCLaZRCG2YlE4Q6tWmS56h8Hi4NRY+wN8PkVeV0rt
zEFS8TTnb7M7QzlB5Gqchv6H2Fgc87+1xYLYZOZbH/Bdr1AjX8wk5Ul2heu8XgE7FPMXRSP0mwE+
RF3BlCy90U1Y6llwYsDyEuHrubt+WNpyeg+cuLCkT/U9l0Vh8dNb2k36P92UmD811V4raa+yucy4
epM6FgB7YJJiN+/qrep1wmalEmMLbvEQcwPi69v3Bd2BEmIv3DOQFvVr0qtx4cVPX4Tkt2R6OcCQ
YFx/nLDMDynUwsUwLD55tNMeM7HfAMvyvTzpI1expa3y4WBzDR7vq45pytIsQFP3WHdfC76vEcJe
m3gaEUCGevJJa18IASfhgkyjJWo/VDgEciNS/ayPePgAxkhLA0iexNMqSQ6NRtklx/KxzQYSTX63
oxnIvbAUAZsDYOmSpl7wlhJecWUKyG/tw0NLwOnM/rGC917aaKI3cBFO/LX90v0iGKJ9FESgvYel
V3ft1IiPtpmna0IuUq6cScTYKyj7CPLRBmasIKVbfrXRtcWppRoOZzRLA6+wWIi86EEeJG2Cfo+L
blFqktGcqn5RZ7AW0l7qbWFICpzXL6CkNiCJoSjTjoZjtzy8gJLVVipg9p3CcivAXM6L3WjS4rG4
x4K3Lhi79DAOpV+PKhPwhGyMvwl8oKL1UqMPvpcCY7oQjcDbLytiN3Rq2uPOdct5EhkMDjaivo6+
HbQX0b0aCPMe0dSJm4x3pavR+oKFEyXszvzJpAK7LIYqVzntX1xdOFOCsJo7gOH+K58ODBBkZjun
BqcO9ZuRIargyRpNwi1qM7W1EHdFowNqDyQK5tmu4BbD/0Is8+rmmfcemFvQ3OzLeFycsonT3jJw
vO0cHcl5aL4s4pLW+2Mm3sj1T7LK4t24lUcMSm8H8jHhigiRSJTkleHgo+QtOnw6+ClRxs8Lraqk
JrpeoDBFY3let4Q3uFDqXFRp8qtncjadtkAmoEYTmRtDeGDTYrQePhiy386QsHs+7XkZzasibk11
+wZlSDBar0Soh5iSiE2NIoLW4iJdNCQU5IFiXDOCj/pBH2mZCoMayAsBPSIdzoDnQOZ4uL1QE1+P
S6dfmlN87ElqaBmaYOJWF84+86ToNZvgAY9iRNB2T65DAkSINjIxPZxxn5wwOs1mjYZDThYHS+ef
a5ciUveakQMmppvVaC5A87kIrI2P2B5HcT/46NIqNKS6hdg1ofXmSc24QQHXt+ICmJjtTZzFAdD8
JErAv80YQ+BzEilREbmHqZszges45979chi+faf9Bcm48foDXa3oj6gIZraI/PcmRgq/nCK2SQKm
cRex2DJGwoISG4K5mrRoggZBLlTqf+UK1r+KXWEXa9XjtWXo9ISqEqmoKc/cIMa6agKja5fkJtkV
xYkGg/cFHQY4ROmDfcVXepsyCkdsScZebjmRaFQUYGFuesoqWTVMVbpYNCvvyDXvTl/FUOuIZMVX
xz+ojngu/6GBuKf+rWsZPnQhNFR0O0GgC3JRVcvTY0lhloW+CQTSRzRCHIqFYcARz9PIEBetKhZz
RHzMt1GiXoEOY5Og2F5Ldx0U7UQsJboKm5lR9yrcZPf6BNRffQKOhfO9Pt7HARs6rrNjrP5r6dqs
sEVMvG7sam5TwT7lpEWFE0rquJzROCW4LJ+if4te3j6DxR07ZtXi3PEQmC+rFzCR02voykJ0+S7f
9kag7Fdf0Be56TP41u2HakzcEBPzBbFDX/dWvmhn7AKExFC52ZVXebStk1RZYe3DHmTLXRGY4udx
oL1hXJVHHEzG3BnbY8RnyLMNSZbsgk8J2Cac9lPP4YlhNllY+lgXHG5+mxzdFNbLPza/VXNovcar
Y4AyqVc/nkvsiaaGa0GqoLqBNAsM/oc1nAi1hZJHY6UXM9SXQc304My3lUf0kmiiFJsJvHvPDoGN
Zhgw1gblBRfphwrvA/Dvqj5d0ET4hom/0jRXYHhyaZtDAdbrqMKPRMI4G4pqH4/Q3ZR+IDY5tGyt
R5NHWl3eclncuFjExnw2n6GYexeZjvqh4pWQ11jDXwmPwUAC8U+wUo8bfxntzGRuHq3wzhu12aQ9
mIzKaVk/POdJ2gRLPiazDC5Nbv5lZr7H+N8ldCkBBJkEHW8S6R8dCmkeKoHh/0+VaezvUGgsCKjk
5BUGi1ZTweavXPoPUx/XLRI7j0smJBPY33Qea5WaRnqvpXAPFFee/wy7X/VMk0cbX0YpHq3Kcesb
AEJmcmqKHTA0q/peKOfXxARuxzPgs9o/ehBCoCWDp3+RXmo9bXuRG+Lw/ANC8XCR0TWqFPPYfcEf
WtxjxRO5GGkvmOeRYPvg+6p0NxMchxXTK0pV8OsECmDYu4qbJ6j6niym8SfHKZKez3sR0KpC24mz
oD+lgwVXyiMwMMcgHhlmNOeK4/3VLQGb90o98JiuSVfr/ix0/YQP0EzoOnJ3L45SMS7fi6tTzQyW
aN7SHN48jcXDYEJo+pxN2clJakt4FjvbPsFdrJLxpoEC/l3ZDSPF+qpxSZE/aTubth9j7O8KtKVv
oqKZRJAi/0/SelWwb2jCFeYnsK5ztp3oQg57SQ6q2ZI8o4TC2CztXi5WVBQhwT36qMh15yFmETKc
Vy5a/O6k/+hH8qIT+9/ooNKTSU8/Ft1uFzdVdMMeN2fEj+b4qSfJKz1lp8IOC2PW6X0WuFH9HS4A
tMvNBi/1y57jvqx/9PhpzRK1Byuzbjx0mLn9gWxiYTSlJcl3jpHj1iF/yxhPycgXA04wfIwx/Y+/
SLlhtYAAlAEZiHwEbD+7pzjPpdoe7zPJ/pz5yKRYTB3OIvNSENsoqHueTZ+5VJIvW1d7ebeC9eP4
VG16GbbVdWc7D5ZtjUTeRgJJOOiJwEZhiMnfAPAfUXDcQF1pf5xrQI2B52sYLV58yH8J76icNxxc
h/tMVzk+9CSKVgqNAaoshH8MX0QABkaD30frDU4a6paKu2Zh8z8URSV3KLvM2TYbJFndxvxv35hG
XTwDDqMUxh8GU6hTV4ZRgwh7TYLb1d8UqDcv0d3LdHkegKotr+5s0PXwOtlp1mOY3W86yv17EYYR
RVR1oBGb1LvEn5zWWUTq+zHLVmycarqU3x68zHvpV9QOQ9w4FYONMFCbxRk94D3FHTjO2AFazK0x
M6CqsbFXR693M8zSffYAQVeADAVu5EXKgwDms5XFrVSAJcvmj1kiRiUDJn3XAkvTG1uevHXV8hps
mZ8fSMBuu5BE4TfPW6Rs1zDxGh1wLaKLN4aQj2HJ/6H9jOfiWYRBBUPfE5+WTnLiWtXK492nsLBw
/XjQ6Va5aPeWGEpV1R/oXFvDYMgsADHTmT0FqAHUm1mkh0jeZ52Lg7aHkHq51ZZtJZpCKZJwLNm4
cjIqGrwUPHOfdNrAUZl3YGD8H4qA3nXrywLcB/1ChTIdcXrmaoRee1mmZDHAGBQ0Bmm8VfRMfl+P
htPkyWGDsYn1aCnkc19iUIcd/8ERh2cWyV4QvVelY7iRytStyo7yifW+mdH6B6MP6nNwpzEqgkDt
Gvga/KlYrY2K9CD38KH7yltOU0PFTQJ+m4pTVpkzjeCyrhHSg9QVaVvjQ82/IalTxRBoJcQaD2FG
gyv1U7CeS/N7Xi+Fmdj2GVZeHsx1lEa7pe1EgK40xUiEmKyBpnhC8xGye4fREmnZ4qf4kPVZzyC2
0qSeaPol4g0l9tEh821OtuSApsN5X7D+Iw2u5oG3MP16xy6xS0t85UQxaPK6YGKgk/PIBr17hDYD
7Q4+IEa7YJRwomp1UVwVF+/QHoNvOKhdhMV8OSsrK1yGpy8XXLpsa2sh/UN16NlG3XF5h2aVurFX
jgEFnuMdHQXc3QvmjIIXTd4EZm3EIHSJxyes7ap/o1CbBDF1DdUZcuJN8KECBJLWQhBltZPwZJvc
r7b4I3hwzd5U7KhXunftv+EMvrL/HKqQVFx2Y1kdgtcyQRAhRxCnAKDWtXPsgKk6+17pR1LaPh53
9ReBS53o5jMtyywv0xXzh0KzkR29GVn2i8uSQLKwo6Zdy3CYHIizVVpn1Bn5Nbe2T1Hr8Q/4fdw8
fd4CW1zm1VSIQIFNeaW7R+jfzCUpBSB/Q1oLjXLhjrJ3ZtTBEsp9PImAx9YI3MEt1yKoscZRbVLe
IVuTUAB/8Wq3rIi0H79lOwMNhsHIbb2fmcuvH2rFihXoTHG89JiRdITZypdENxD9pG5u7hkICb7K
vZyl7sch0Z0ZcWgz2CNJ8BYpyp5iIJMhjxVD6w+XJeSBsrWbEqsNRdrhhbcJnmSBAzq62R7u+s4p
iOFDbaHwhBl1o7oT3w02oX2Kixe7HRenmnvjvvSkr+KFWoW0obzFJxnV/ySjDkdCfURjDlfHHgL/
xJbXnnM0XofDprL+MIkrjR+0ABdM/CKRkY4OBVfGxNjqs/NXuLksVv+IEBmNXeWib/6mwO3tpR0x
xWFL3dSU1tGARTehnfXaBkIZ33xdc9YCtQi6wqQgDVG1/u5vLwPcIVeVmRXu7w1Dkc1Mt3MVs0Om
q5zY8Ju747cZAOUDTK37gqtiyQ1N2Fd7FhcZXOEBE94M3+6hR0qJ6GU/64sxf3M3H780i6Gdr4yM
2QnV029hLLZhD791wz6Wsml+4SQIgdSqsz1V2qvi/crQ5kszyq7fCab/gGYTNnnwk97XfkHfrj31
Wa/BROTtsuLTfC0JeocX0678wA+YL3O/11VdYiELvcDYXuvcnuvYzuKf2X1Pj49JzW4zxS0bfUMs
V+kXECqjskqEVeexRNvdmaaXcMruBOxg6VAFkvwcxLxZChlwRABknoTh6OWATXsWD7d9ibX0ZnZ6
fky8fNIvr2wumrsH5TQgFKd+z2S9P9zTWdr2cc2atd5SyEy0TjtG6r6oaW5Yhh8lk72WL6TyZaDO
apY2m8Ur7O3CRFo7kXW1NQNCc42W7U7ya+ccLNgtqTpRjKqhjlFJQvo6zZfMVZ73y73lBj9eXANA
nhLjWSCb0eNILhPCkEbd9jsKeGdJqzmjXyVyKdfbWQOGqAmunWIChTK6X4zIFUKxmqky8+yOSWXp
vqx60EoGYCf6KuhGF61bUxX/O+pfQhnjrBq05bdMUeSLmzsgZHdATHMjXawAO1OFzfe3fmA5CQ7H
iaRckyVibS2H3jX0sJ/inNem0+f5tvaqIgM7nyOGADElfW//t8019kOdCx30CwD6LTl+Bx/LQD/1
DlGiglJJURBsnxvVChK9o9XtmUlXzLp/s9COLwARHyedsWxsTID28J1ktLDXf8MKXaAfU8bYSGpe
NwwsFnzaKtiJ9Ww86JVWXSKltKgVQlKylDKrGEXb83YaO2KOFqQJURekpSwq0zFaCawWXrDJAU3/
/lRJYPykt0wOhtyNzGBKiK9+I+ClOD9jlUcTTlwc+TIhljxA1cOY3jZcTI3hbbMlorKtBgVu0Bqp
CUI7foCVa5VnhWYl0R5ROv1yla+MIjkvYvBIZ7c8thymDlEaS1qta2BhAZdr0jr5mPoxpmBlZB86
vqFgdw9Lo/T54SHmByNrR4Y3cLaCadMBi6HdrkBnY80Y9v08h5FLXSo+VhU17qovWuRTK4OASBkr
Ld0ZhLo3lBa164Cz2XZQaX39u8aIbJL1xlV0urO/Uy29PzemqwbQZL8l+YoM6D/L7JxcMkT9rzFQ
gI2qgjXhK51OGKGCSFrVFgBpA1THtN0DwF6BkHdsJuKLX/ovGGYRG9fJpJwdrlRScLIBx/PqJ/tm
JmA0IPeIpEthC49W/njnU3d6tJOH4h4xxhSDNJHvv54uClZxUbGrDgpJDaNLVjmK2h+Q/VRhcbtB
BobfYvh0WSycSlo6uIRimBDbV98sP+xAYPSkP9Nq1oJMd07hYc14OpE1b5bg4XpksTW0Kxl8CF+O
+SQWropxPQxDYwr6JLBQevltFdmwzYwIEm038zUXN5Dl2KSpa0ROYa2mguiFnX0ev5m42od4Ich7
hKVkvmviQcV3wbSp5e3ch/hWziCVJrKtqHGLN/dete4o+AiCaeqlShWDz7eErkWDR5z3hNfC5EHs
qwRvYe+tVR2oucIB+Re2pud5YA8iz/pkaLxm2Rdz0rHIyo7bgRbdgR5JWK7jnj9Jb0Ckgy3IeRJs
o/rSSUOPLB1hfN5kDum0/dM/ywblBEoup+6pV7LE3t6/1vgKQFpqZQ5/HLEEL37IXzxRxV/ecx4I
dyiC8vtmoJHE7Jj+Kf7z1M3n+9pyiKcvqQvDn9rpwdAn7L6UNNEuI9sKg2qXGWiQrO6bVdqfyodY
elp/5PalSVoZh4uK8GdY2+YEWboZX3bNVJ9RmH1pk0vSA+hPamiHZq1c5nasOyjgPlXuHgd4HNO+
ewVHdpEFpWlKawMm5P60VMWIZpDBYfMFbzPp2w4qzCw8ADUHHLukSlLaNeQckzydNtSLxuFADO7g
WsOF+SBN3BcbwduzundaLJ3ce6TW4I702DUTBbjsV6IGQNG1qTitAMUE1VIFwW/iL++0jEOB4+Dl
s1+lxua3X+yFfe6K1whMQ0Jm5U1Nn1zs8fDo2pMax2Wt3r8TKfCB4nk9vmhu2f9H+X2DbGSYWYy5
lNvPwDF5k0pil1AwJRuoLPIIKWt4rHOwG8FgAJbfLsDZhwO4Hc+GBJjLrwZTzD3sCIQZrKP5lULu
Ba8k44nBxWemIFJ/z7UiGqDAqEZEKd/N61tTtko2Cpx5BTPcRTioiN4cZKLQUECk07iXLWf72E/V
R3wALUlS7DVzT4lxSFUjYydBo+Cbon+rmIYhJqLMsYgPS/6XrwQlfpe4Cv3DIVFA+9EZruCKPGFJ
N14P9jNQiRLQGUlpbgcoN+1FzFD1IyqbUYvhSodP3GAkPUv3kd/N2/iMvOELdrjPjOMFSq0p/2O1
PSb5exxGlwgNx3p2OsZBhsn0mlcmfJn8AVuzUzlSei5J3Xk81Ls4huqwHJTlhlUdVJoWF7CwwNP9
tXIDnIl3EoLPVZp6fyXMb0sBO0nEvaf9a9TpV6y5k+F3KL09lWAQwWFqqUddM6dNa620lE1XcnRs
Cyeblcrnldwq1D8oqgLpj8g2EB/Rx1VRooJA6oG0ew5MgGGw0b8EGWNWhNmCsPcpcLSfm0AIhlCF
m9q6zg9gp8neFNivMPBMznVBern2L2TkMnBI03clmd1+OsNDGWvCuB/jIRp52rdCh3/8Vktgp097
q1OPRNJ0dsAIK/1DIiJDlnaftJZBlo7GKWf2WMKnRN42utQHA/lGXOvFME+I0gloyLdupCn0cpmk
havTPU1EwWyg8rnizdEqykcQAhXaJmXJPUE1RPDf0xAiAHBckKspEsJkPJ7DCurNvD8BBPCGo/ZW
HX6jlhvVO2a8+7n+NzVXyS4/kN0PAGc4p9LG20+3d4X0lrGl5JeiRPsHTNO8/kcLFxiTgKKOUtpw
cSMBHLcArgtChHLI2zilL67Y72s3dmrnEZ0D5znDxbYMtXSuvFdzl/Nk0o5aIwIYHSkFgccFZDkC
w3UH1SQNsreWat8eslA27dPEYPpJaNV+7GFxwd2Fs/7kV/kMHI709MxGSTcMsvy5pxfb5comtCrg
F+ruGcehKgoyA4OC9FpRUDAM8ISRR0L6+WPUIO/+3N8A3K52i+Ea1/XmTxKwku4i3Tnwmm7P9JdN
aFf/fCCvxvHeNYdeYxS6ttaDDZ+Q/kgQxr2HjMqc7zxCxm8wjnZMOWSoAjfbxUHMMuV9phAS/pEH
VQMstrwbTqaJ2AfcVMNRPXmQe4KA2T6nyge0UGzkSy4E6inP+SHKyfeD9V6KnwYSGVKBh0IYAFO2
cIJFnsIqtxSxcXU938/LDFN/iMXgXdFC8d3d3CB7Vu/M5QI8lAYUriTE5GJf4lyUo5xdDK/LaEko
PnJEk8ii8qM6ZsY7xL7+8yczjKYFotXfSD2C4WSbjgiPOA4vj/Co0fubBtQ6do55/IIj3vaeBi3Z
q4PA7rJQPo8Y933p00o6oKrrt/B1JzLNYlkp5GoVt+eEa89d04nZ7ync+OaD55lat4rUGHc6b24t
X+6bEZ6MMzGgvj3Ow8YhZYUOaMkxiAWnuTMRIt9ahUQ9qE2SRDbrciQsg1UjhLjXe6wRdAOX4wwa
iu9RjlGq1/weXFN4Ka8SruAzP599YN/RMcg3p9TvqMpGmoyo6pWlxC0ilzIbDTLblq2Gq17usesZ
O273ESelBBWsBj5O6ntjcZ3bwrBGTXrTGET3IV1VrWapMQkDEdeGIwb43hZBIDKz2hw+ABNExQdH
bqOvo/gTrl3liPYl49MvzA5tU0+XM2dlf2a9Y/VOpTDZ433+Zf4maR6rqgd58xp4qeoEK9V6w2GY
MTww6cB13ODvFUKHvNdUsxairH7eCGJgwAyOQiRSzYIG/oPGoL0IUpiIHoxn4ty43HqBg2fmHasr
iHbLMIiAHKc4NzQKGFYT00EtODczNjh4Q3Gap5j9LOm7gkkwDZc1hWg7tjsLZNZCndUoJM0QtD5n
28BfaB5jqi5uZWDnIY/Y3OQyr+U8NhM0VHgZGSbLBaBrFoz+2Dsd21t5x0go/YMQ8HLUcCDaN+c+
pAokfNzc3WGgEGK8pFwQu4bd7arJf42hfS9fxjncXjPkoE20/Uwsfzqz52cbnIENPZ1Y7wj7kqw7
+fs0urqlpbGtfCDDrvMsKLhZeBqE0iSKhnhicjUKHoL6Xu/zJgCNKY1MCm5JIPl4xCXKg6GmvSZS
FQml9VICTVnNFAN8rOgjSPpZEnLCKwdZLrBi8m+1xwPszwrwfVzZX7bQ1z9dnIw6reaKttMA8Ftv
e2Y+JLvHTiUpQ9QDxqnFEL1+7oLrGLQiAjFvy/vDzTscLr/MlWanYHbalO2ssV63G+d5N4lJgtXA
akFIy21iZOrPawJFFgDGj8jvk/rwLKM0yOKqWYPzRCu97SbBcFsJKt+lNj/ovDu2RZbydzXgLzhF
XoGxlNslyraRxrwKAcekNrhQaZV6vmxKreZ1irH9svxqH1BAZLQGjRMsIAiVxOJ34/wzqlw26Ly+
SxfNJ1FF1S2iEHjr5+nwbjYBOWS0tHyzRTr1+BhJyrEc4JTDyYI/sN/J0irJjHT8c33Sl9NpnL+a
scp6sIsXf6v016dtPFW5EdTjoXVOkCVOb0R3/U+PxuVl/cExpNMmAW7YBx9XwY7sobd7cyMRObLN
aFysia5ZSqb5BnWJcTVxS/rhMw1vO6RlkthBK+ly1YOd8ZwwFvebyQP2zWwvZRhlkgcertDgNum/
ExAPuEW+KVekYjh6VIwsElVr92OHrttwpLLUEKdNHdd882MMVGLRhAYh2axhGLhmOV7kp5A/vj7I
mpyI6eqaDLblc4asWTmiGRKHWZGxuiU1e9gdu5YE4CSgdoTOHKKC0Vr8vZ676LLGnG1w+VTXALjI
GD3F1ScSL16FhgdRe+umtWRX9Qj34s9sMqueVy/7hEwelw1y/8y4tN0Gy55ZJlCQ+wLA0oJPh24t
rlCwC/8HeYFRikm60dnDYheHOq3UaNhJhMZsTUcKS5Kx6lFbtiRxiPuniIHhgKcBHFCCs42YCn3B
5n4h8UP7ZWe9uooIVpUXbZFrNXpEzy7LHg0Q1dWzq9IQjYIzYlY28ilILoRL6gXg3QXJJR7ZdjEu
3nycJ8jeWwLksuW6J8JdXoAWZ1ngrQUeUVnyZO6QnaKjqgL7H+kvNxIeqeetC697UCS/SOk/Nqez
pmioWbc3fY+yooPmyGyzAiAaeAC69HeRHCS70Osdxx7P15qoJ0HWNy+n2f6Wp5ANN9Uzxz1sLqXt
iv+Hi9ZwHcQeblx6w0C/6jLjR1f1nrxmMlrQQ30x0Wgg2uQkvcI6MBryD4cxhOMwmMsshJJt2E9/
UarpAsKK1HWeaA9RQNG/Mp3KwEkhVYIZZInuvpvB0LOH+mzhEje+0/sfb3fQ5n9pcI/RLgXCWXtO
Ygc0fat4u4rB5Puh2KnOrAAbbXSaSvJgViIuyNnYzVNov6Mge86vB3PVSRqChtHMHL4uxe1t7uL5
4975PMAXC+wTolO4IEDMU5MtexOtU4vgMzRX0TuLL86Hp9PkBg/dyWODE3yhTSQoSvvUSIwZgg5q
bkeX1Dbt19mRnYWvuM8CiwMCGvdu3vq62ra0vDjjemSnS7sJoxtxbJiiAa00ELNhAzWiP7j0CVJS
Sj1GJCgKypTaUFprVRIUBEcNvAgRrcKNVrM64jc+SYXjTVxer0N09uNjA1Qk8ECtP8gvMpR2ELYb
liV4auONd+0pKeTP2IjmNtz+zpupFyMD10EgEkG80Pgqp18RIpYgajIxc7wiv2orJAAuvL59C6Z0
lX07axHGAElRb6lyNVyfCAXa+JUpYQn7XYw8f9btcQ/D+8vLxn4uWjyI1DllJJxqK8E5gwwZK6Qn
fJHmqmFHX6He2cmnk3v1F26OoEJhi/l09HCtAAEGDrv3RdaKuY040yyP4jxU3BMaXDKvdMEoKhww
4oypHJ+jWWk88xu1/Aq7Fku/ek+aOmKIHDUXrgJMobPbllk+2FtJ2JHag6NK5x6zB3gxxQ5pVpPB
svN3KMWi09ZtaU3t0vHe7SfU/BB16EVy0CiGMew0UKQ0uL4OkWa+jMpATe7GSDnYQ7IE/MCPMK/M
+XOQ3G0i6XhpR/Dkl6TKHjgssdrsNr/mMEncfK2Upa1V59AvH+5B3ElVxBLCOY3diHx8o6oy1Qel
cdaqVBaS6DnMTb/KzlxVBzxVtQTMkVBegjfuchHuhM6U8aE9M56GpVnz42QWHvwQMPXjOpxC4PQS
T4NaUKl9RvYaWZEdENgSCGp/P8zp6NUkO+1smAdrLUXMpuhSVZrTAgipCjTvXZOW421CpkGB6XDO
Esci+LRG61ZbzvGu5bOWlLs2SPmgdZkJYHsiJUQHoFg6GKTXd9t+v37oOxzxRfanmVKEgJ1Gvd+s
tyKj8BmM6n7vHAal+SNw3WYFqkW/dGWlRdwyhXGWoZ4Iu99tWeK2dxbVHbJMMF6NO5bODeZoh5Z0
GbQL+hmtjw90EFE1ITyT5aj8gjF9u9CH8Q6J0SX5m2/c/MVAwtX94XWi8ZJDiQt23hdc9LD2vfz/
Zldtn2FOdfijbaQzygRqL6yYvAwzlQzcXveLEhInS/Qy6UOtJEvHqXpClE46qBbPca7ygl9H4Ztm
o3AMNWzHwq8zp5/45tfGWYf8XCpiu+jRi8mct/cWnOpyoNKiL9aPfUQNTNdgK2cq7XqrSKvZ7wTr
LrhffAWGz/2ebFBYLRyVNFb3d9KZ6R3RHOmZnGgJxbYXS0ajEAY7oAi46whlbtUkEUZhGTydlrtP
ttvw7QM+CDJEwm0DbLbVJ+6b3heLmpRTwGQP1VOux9IMDRCFl16UZmu4zoZzuicCqzBgJ/kXbR3b
vs/Mlt2zt9hDV8Zym5XmHFKu12xaR39BX8EcZWUXhM7D0+9XLwHLCtueSZcld9Xd+C58okOxm9M8
FbEfbq1wFQg2PKmmIoeFMR4u7/MvO5J6nuYViYTHJhiqIktrsduvM+NJmqBA7nROgKWCp3Kkhiiq
usROyY98Iw/QkXNFzIwpvEZ12o3wJapKNj1lJoaHBfgNQ9gYsgl9SoQ+UvwRNNjb2CXoUV22KP/z
4ayu4PUUxrWVWuelGiHjZu7Rot4Tvqo+VRCKc+cp8dOCilBfs8JNtS9DZ2WKCTNWeYh5YNPl+yLk
2DkEq0QuiLwwDe/KlXS/b+kEodJ3Z4FRG+ZP+P5qwnAYIeFFhXJxoaRPme0sMhdLLS9E5+mdoD2M
A41EJug0JQ518V2EmbNW3dBkwz3PnHmdIBecSZmQY1ZrSEaq3txeiQJPr7VwMDgyWq7oCpxT4q1e
P/u8E2/fCyWXFzDGPkVsgaeW67QgZoATJ41J5jjt6iHQFZtzotrOJvuR9u+cBYlNEa1Es5j9kenP
5EA8YmvrUhTbduIt5cghGjfHpr9lLzIimyqOk8vKh6f/O0zZl8r6e4SfmzVW7czIucWkuKEW1c8A
G/l3zUiXna4YaF8T5YIoOfo7/ETXCKOeYa387bFb2xAHjMGjdqr3OEJtmpW+J5lahNw4NpYiHLaW
uEnZPd95aoSYgksbwMkSfedmVcte5END4SunS/IwESblvoWz6J8U+F52uHokSb7lJNQZ4mzrGlaO
OxnS/HstWPwdGAnEE273v7YyDzTGv5YD2fit/IlGYjvTEBJ0nw7AShsTmARNsya1qCs46KZBwT1Y
WbcO6h0EM5QGDrFP1yKjE9xcOzwGhZlztzIhERi7BmOZkt0uiElVzq7Y4ADqEk5ysjs7EVWbJ7Ox
V8gtvBDJ+bkpUZnyJw5mlTtb/NVbw78/XL4F6dEq44mXZedEcfdCLrTMbygGR5ZcOvUnnwDgGNaA
bWQpSGh/uAQIHXBPB9baGp45b4Iuo2234veXtQZZvU9zfME/qtN9Jo5EXHxtICDzWCewUF7YXzjG
eePXaX9hwyKiPrxkX0UztjbdXrcxKrPUaoTdq0eqERuECegS0w5vzFhTC0WYpTPrRm3K8AwEs+3X
cMU0fmbFVjAIqILB7087+y46csFDkdlrG312v3U05mMEzsfRZm0mR9ob3fWTCmKocjZ4G/Nzj7+x
oGZ2sjRoXTtQbPJzoWbss1SKGAffi+TLUujdQEmPYxpq78jeIy9GGC1DceyH5Ynt63KFZEMqGSLj
xmpjqBDaoHxdKw33Gk3gW3geKhXSML40411sB4MfY5F8S1JWB/Iyh/phK3mmVmDDKB8xK85Zlq6h
jP+Xucs3RilyhwbUBBZWDaDioBo6xMIMUYdvF2lWKGFeFQEhe5cFGpKwYkxXjECVUW8yQ25MLkkA
SykufveJt38pgf6kuLI+fiOur2yt56TBBHRO3bUnlLC/PyehRxGNI7JkdIy1RaUzs+A+vACUkSUp
pWWkLljVBMfiJ6Wj6HcdltDn1NuRTH1bQb2UDdg+agSl2EMqhHqAnsb3443McZMFjfGuoM60qiCK
xHLMizXviQ5uW1jTTK2K+s9z/G5FFM4AgC/k+229zcnOzC7cE1/+2D2YO7uwje5HET6tWOTmYOv5
+XsDWkk0qx22xWHpJqvtLrYm3kfm820uPkd/o98Zrs7MXawf59pSSgSXAiX3as9HSnVxW0Dk53Ms
4sLfwjr9GcdqpJtp2yt+Ni9vH3o4p+v2KZdoGlkUsjrRkECuKrDJCZTTQ3i0mAabY3MyTKMDmgji
KeIBoP8MHoEx4rQlk+t+l42XE8/S86GH+Phw1sii7dkR+BbnE+Wyrd2TX5bJM7zLhvKJRfcZ+/Y7
YUcLZy/4xSqt/VpIRONSGfk0RGG3GrI/ZfBHCUs1WQxuctdChf8KOYnfRhTWH5nZ4+9Y8P8YA4Jf
mIkEkROTI8AOCBspfVmUa+ffhlqs2yJgVnA8uctdCc3wosz34EUiYTQxSH2rjofyOOgICXQvYjjT
gQsPGRRDQGmzKYGt38Fr0FwyyYR19PiV5pHquE19/eoL0DyMMUs6+BwspO3bsdiiaglKVLyAS9LT
h04iHaQ8mHfH3xUt5kh4x2XmXNldUJx5lEUPTqFupWx+HJqTQ91arz0zQVW+4vU9l6znPRNQNkDN
rspiUtxL7pCmBHip6rDMfuIe0kfePX9xEILuGN4Q2IFPQExTE+kHQeYuxniivWwUCs9EvNm7XpsY
ooMKS4v0DLWzOReAFny2odjEDmjac+AgtkcAwEeFd7Vl6XAb5VVzVoOG3qDZ1IgWmQ5POcVeF+T8
AtUWIu0ZWUkskiK2qKNh6Qa3nZUs+U+BTexHSlzKyjRWpUSVo+y+/lCt1iJtaowh/HcZJaFbu68m
Oex8I1x3oOg4ldgSafOcfGH38svNivs/rbUNAvkAlHGdU+NPJVoGjcRBhx+Pk9DNq8Bu9Okfutvu
K55t8yfj3ykb7y+d99vn2JWUQbz2IKwVZ0+/iShMwpVcf2w+deTSymhuPml1/Sleou2omPTzFdWO
sOkt6Y+5/r2/OcJgs4H4kTBjgfjbIUSh3G6EFd27QpWihs/8bMwZRDzG/brbFekpoYTjtnuhG1/+
K8i9K9dpGsEABCd9lBGLJpJDtlx7rRY1hufmXK7q+UpRDXb6oSHU7rfzQem5UgmxJbCXe/kTpf4l
zLoh4VSPhlHIAWsVQmZWsLFoIpe+c9zGHR9Gva4MguDjyglTezn+iYwrLVSYyXWPwgj7EmDSPIkR
Bzt/lKkO5sufN7J/c4X4KVD2m6en0j0ewaAwlKgJIRAYK5Ein2AvwMFGi1+b3EESqPF/HuiRk4wn
fXon7JBVuINmJrEeB526Kz0eqfAJncBVdCO1xeKm0SeqXjpjSTg6MItvIu/c3yBuqFFYtz8wmzfO
h8amFtGqNrgMGa8CxzCY7C/lYPrgLy7RJZY8J8xt1NAE9kDjB1KOCymxV73AYilyY/KvMLUMuFbK
Yj237TbXxZLHHYptkNPQhhffbx2fdrWnE1EY8RmXlyLANvLSi2tC/iytblN4m67JRKZ7s7kbN0ug
9XDXCADxCQfP0woZUqNZLMg2olSYR7TlL7QlvmWI2+6Twv27A8wDvBIFrBqpWwZuer0ou+0hGhlt
m3EzPEJ2TL3XeDhKzSmoI34TUvXOnyjsMk92znh11UMfqtAZomrGOrFjuJGxctoSY3RH0rTBpDLD
8XwpldUy46qm0AC+6f3ugNwHxtmWqrRcUI45bIRf1QB1CnYt3fcQ099TOSHmCQDlvyV2mnHDMRdc
BYwr4I/c+6+ai9qljggUjonjFNIqrThBjIrGSMt0s+eICqPjV1cZnqCpAzoBG9dD4JHwUUUogJPm
GbQ1+5s98VBNBC/yedpZOEdExRGDrULCL7wEcDd99Le6A9nYfCWMWXQG9mKKjHYy36J/ai9+6h4u
o7bzkNI1wtiYwyhUXmSuQD80GQVIvS5pA2MRxNoFWg3VeMKkVoJ5T1WIsJh9r0QoT2QQdnBwyRUb
4F37SU4azSuPQyewO6VWTwcrHCFzr018h8J7K29GR3rMYk0oUAhdk5UiCWUj/Y1/nocOSkirfgwO
/dsZq+6Sc7hAXYWnHEM4eBaBhQNwV9QR23PCFK9ln+v6wOSQUcvEkTyFUxx/KBPgPHnIOTyHNdZM
69/dhKSz3BBzpc8XVphRNTJ6pwxQcgAfg+ZgB9uGmZxWvJxhj2GgjMyBVp78EXuMAtOOa7XS2iL8
gPC4IuV9g96pvm8ontSfzhk/LUkw9M0LBrftTGGcaBXmRqOSxbizDT9QkaAq9C5O7uHo/BGPfQl3
oTxT8n7ocgAuIcuE9xi9CwXIoxm2pdAw7VlUd8Rnc2rAMCf5DgWiTuwAjKcSLNzJRuxFXEk3So6O
RSEfiBaAEtRpPU56U6rEFevOzEAb7/nyhoYiihWDBEpvNy2dy7pz3Yai0avdg760Lr+X9jTFl2KI
E11DktAzYAQyk7jgDzI62Zm6uSFPo3RCCXdkcwUYuPIsVfZmmbpk6qKXl8sKpD0ijTmQNTvOwJaB
QxRX1vKWl/Ob9FAD8w9GajcajStfTLeb8y+JzwjFQGfkcF7HgK/O0S0SrzJfcCB0mZyrCC9ZevtP
c4dqxh4Xdt886KhX1Am0MT3s+4P/v/lE5WGwVZaem1+Gyq5MPnfVTp4uUaivOdgUzWdxj9u60Sr2
+Tm9TDczeahfjhywE23YyTIIRAOE5jVuevYPY58bFef3UWNSic3J5VHsrB9BqVXI5kKNXx/ZU9vu
xXQMwA1ss5eyrwoJUokrzKBBjCXctGSiK13R2OJ4kBoHOIjTAoh9DJb6RFf228+n3L8/XtybxWhm
3AChtGFVNh/tFp0SIZOy5E1U4mU7O7Qnp97cEVKB9n2nQZDHimtGPzTY3ZYaXDosTEaUjsnonCOo
K49+c2rnfyOlJeKrByEuKE22yFlNcQijlhD1rfsBliOPyec4/0KA/AJNCS46VYg3q6kwjhZjtLRC
fgJ0zP5wcaqwPbtFNhX9qqg7j1fkkYWMo+oaKl6zSyUXefAIGoYKkK9RRvAc+DlwO8KQ0sOwNVuj
VQPnXWVLrp2AU+7n6SkyeCO6w7sMPCxhD2O31VaVvSBZn8srgfmX2+hgIlkPS0ht7qNn3SxcWdkL
s3UF0BCVJ9SseL/SpXTpaCdUhww/u7uVVEIdgyyJiCPQL8W/fB2Tlw5vMgH3N9XqwvRFK7f0jEwZ
xBlVZxSGaaYA2Zj1xYXEA2CjArKoUQemAn3acxmjvTrmg05uyRiobdjSp4HTp2vbzdkE+N5qniUo
N8m3r6QtajTqYI2bXGfXHtxUEYgYQX3tXQm+GIaEjJKwwTv5zRNEuWwA0IOyZj+rL35xgZpr8NCe
3UKdsHhfQOCDCpuOUu3MAYtloWHItVeu5Q/g4s9LwibnRisESYWG6sSzd2jflYMagnGTMNsqtKNC
iS4gZYPqpOeioZdFY/IUTGDyEU1sQdbcbph7DOztbkRa18xsSbo0KrG0DChc8peMLwjEppFnu+jU
DplU9taLZDvweYE0HHdteOrPAPHp0fUg3v9kwPZk7X94IBhtv1eh8or/Ghp9kjYsnxvUsEL/ZNYt
wY91gUbOyerqM/iKoAi12akKM2X+h61YHY61V4bf+2QQyRrGFyvFJspgBFYXMHvnb9epJwxh/yhw
MumTJnnY6PGqeXfYUxcfq7M6/xrTtMzdAJDesGHd0ibYENa7wouThUuryfny4YXtAqATiDB1Sspw
KOe2ArWP1V+beU6ghJqoRJvfH9XfOXwlSAsYXmpRYg/uCEFK5mxIEiCxKXxs8VV1DWJ8HTge8/UZ
XdSjqBEjQInQx3zMiOPTgmQRfHShAw0Ji8ioLvdFDS4b1dVAazuocZqPuLt4XPgysCXitSwzm3im
yqF+9MsAf9ZMBoV2K7gw81M9oZgev3PJ2zjnVN1EIqUIkZnjaZbDjYiVJth/rCaUxFCK4OCxhEMF
rby/d5lcsGWw7KUHPezqtgvHFrJzbN2wMNFwMKc1LBETtYhCmuFmkfrn9Epko4dww8q9xAil+qjJ
ZTcEHwmkI69Nk8/HSdwTgO/Z21rPZkTMpoZfcOzHKAVQEcGJ5luwCI4nHxEhq9VynHRMx0ZxBPWx
9zKPtTD5Q9LwejqT8/Bql0sj0by6SY2xWRiaGpjlFr9G6srrazsGa+eQK07Tt65eS/oV+2jcaTW6
SJFmBFDrQUG6aGByMCe9Z8Nw9BnJM5KMKZLjUtkRP+KfC9LCrlo8209NSw1Uia5KfFZTEr8a5kDD
7lZ1FwVPL5Dfz58N/f016dJFiRBvyArfNrjt4uiee8WmlS+9xiAeK/VGuUIVL00wUt76poZRGsvA
TZxLIRdtt8w3ChPo9YQqEBG1Y/CWuEab5HVB1dyeqvtCeo1rC0p+/qW+6gWi3ewTudgyf37/wnR/
qHU7pkZ0pDAwiDjf42E42ozptGKPtcmgqdu2r/7Ht5MjBivF3o+TJj9aB1h4ah7guNjFUiVYvIqe
kf7ZDG0B0Z83UT1MPWvj4VhPa41fZbaiI297zOkyBNjAh30ASzGrd6cC6jJvZMWgtvcSYbN29lkM
18zJqQnlcvHXx5R1E0y/2tjjbfJFmCduRsiVdueNE0Jn+QLUwP/0SakhXEUVT6Qx6h8oRtQQoQJF
9j+weUVkELNxIljY6svgR+rOlgNcvAN902F7jCOG7WZgXWKqQ/UVkvXqqWvruBto2FAhicw+TDOv
9cCL7OdYwh3DhC6KStn6nWfMgz28amw+kzKMIFPbGTvNsCHLdpASVIL7jKMGTkZluiclmNVcHMyc
ci+G2SCT6VOwE5nYB9RusQOYNHH2LSi4MGvoflLeEa4rcXANa/3f/JCFw7+eqgo5BCHwNo1hvHCe
sqgXyTGpIpHL6rxCGn+ka2ENHIe7doy74eU+wJBip4qBhyCRtBIYI2slhDdOHLDl4KZwLtK58IiR
VrOrpxFSZqFrPxtNzYfFpplC1m+o4444/kPTj2IMwlNYX63zgRQu3UVaAUROgp6dFY8c5IxzKyGL
1WUvglCzHtoMHZn4RkP8Bg3ZZZPbw+shAcNIJZuOrpsDbQ82jN8a90QJ6OvaQzqTfoQIylxa5mv0
Di9+4revS6PMoTDpo4G3/JYOqOev5uiBEvNQMe9FtAM5qXSpFmBToA0krpDVm305mzZnYrXmMSky
jzcZ+tg7MBWohUrFwc7iXDDZ3CtAa61lBsH+WhSuW2p0hh1B/me6BhJsybUA8Dd8iEUTGJZyRGzZ
oA7jA0FLrJWlAo0me/JlYVkgS5mPT8IGR5cKAyEbAyEsGEdxzuuOed5g9IbKeeTGcawDHujjAORX
EbYoAzQGTLVtHXyR+HT0e9i36O/zKq+S0mlLy+gPSpSwyUdRshtOylGgmMsTngX7/yAhm4RM2waZ
feXruAFgXjeAn+hJbTywi84UeRiJHoW/f5r+D7tVOW/K7haK/CqHkwVHlne/eeco4QvgvWdSuCdv
oSQkJgeUyAVUpF9yZYlV0npolNxC+2WA84LZ4X9v/EkVhBinguQMhAux4AbxAcmuDJW6FATURrm2
JPnpD2hPsLa7LEe4U8amci9qBQ7GZWkAtxw7geIWtf7Us4BiFgMXbuxuaRyEEWS0P4fKS/G0VIYD
OwY2ZB8Nuz6/8rVogorQWyAL73zwC43Erj+Xhnb6BS64PQ6L2sMzJLxojUm0RIqZgQlbjlpeOK+x
Sc1xt+x/4U8Le+8wKHtWmCmagD6efjCUi9++3XcCnURDLlp+HS72sYyHunq88VUruwu6rTEItd0w
WzTdCDmbaMB8PYB/dWjDmh6UwkmPsaRS9KMAjrE6azK2EXdAg/x7cPM+EoBtXwVG86EwSJxkWQm4
TLlOCxW6F+SXkV5S6mdC5xQ5l/j5roQy420wZ0BN8AJ97wzOBISvOkFNP5f/ke5UbOQFGB9Ozi71
3iPGSbuBwtS0wKuW9rs4lVlFcLlPYvIcuv+czRILbVlhJyJTnuAXqvV2QqF2WR68k+Q6tftg7l6/
edC/c4qUdrOAVwq0vluaL8O6xoa87hbFhkDYUIIO2sdjtkM+bFIVDwXxsnKFO/zbxEOOHaW2v15a
FGhtaqHvOFSZIkJpSb2LuuhDyKn5CPs9mSvlSXqu92wIbKwGUEQgU+FbZJ91PNhMNKwv6sFSdoFI
U5apf0ROszeSbIeJr+vqS7Wkzie9Q1ANlrglILLQB85/lz6Iv7yir2BD/mPU9oe2IwCmWGOofN7S
QIFznKqHe2oLgAe+ahNtHUTvvLsOi07OP9VfJpfgsGb03Q4pBTVelljzFGGfdPGjQntx0sRR1SmA
HmJfg0FJ5VJaSLXVlamnzBzeWoAZOkn5hhtOPSpKgFxZVQwm0o4doWTDT05NwHtIN5MRc/1t5wys
Ym1569Q2oc8ego3GOaGsl3jupUYND5+ODaJwWC9fwxtrjxps7mBB2140Cf04FnH8BwhYJjBtwU5/
q4E8E8xUth4TSIsLe+7SNWarcrD7JrU8786laYv/aZ4jHncj03V7HsXitrBV1FqM24mo32Yd0Zg8
zgrkiMfJKXmU1ERDf2RpDToSz482iNh7VPOwsuygQmgOiEjJCvEDTk7DJBz6ri9mQK1H0nPbVRhP
CrBKRapvWMYlA72RjrevMmTvyerNnbnldYZRvV9Co8fG50khAA0Qee2/97kPNL5S8s7YH8mLXpOo
cXzAcq81p5uunSJbXV4gnNASkbq4tUlgARqZ17JK8wkK6s3Ctfp0Rg55wBlwOvWrSQsRv/SAYYsW
6tQTnVt9Z+9pqXFVlEufj/Ta/LZqG8B1QFTN/siNTFCqWIpE6ebfu6NJeXkf8fvd1iJHVVN5Px1t
T2nMctfofrMoz9lBy5niiPGQO0DAETGjy2lbXZlYDh0CeFV5Q1e78F8FmC1MX6qen0v32iJkTp45
sjri3f3fZ4q8CdvPuAPB6FD2u05w+kTG2TEgv1/sMPGarHwDUueM4SXzv1HyKYgnXLXRJkGmTFNX
/VVzwQUq1dq0ytfx4ESg9YtHC1CvzKn+zmoIe8hJ1Ub8wz111FP77GpwK8qzeIBbnFqWl0/Kiy2U
BOUNccDEimox0fv2B/aci79xZ/uQkDYZCgQB22JiKtZQM+KF5qDIk2jk1MDbmn43v7TKWnv4VuZn
v0nzcwvF97qy9Q7nhq1ymnie+0dvO0U0Y+sM3cqZ2RY7WUts+t0gOWvHHb5KMJlbgpg+rCnpC8fw
6np1Ik0V7EYlcj+KhSoyJ21oKwGx3i1HwuH/JMfV1XNio7QUEwRleR3Lb5DTd092Cp069P2AAUIn
/5KeaMEzHTG7gcgzpxKWvX5cPf8/daLcaoUB9NebT7lyH+sG2ejg614RoHhxwlurez018uxzB86F
iqDme5JgjP1eYBbVwGcupe+y6pm7rUPGqwvCi/atJ2LEynLegyJIKh5IxtKvB6ZBXpPhxH1ZyHaY
gaZMNBStRH4M2URh8WQjauQDc4yeJky90wtieC6kcMqihm/w0SfViVXMuRXyYxC3WQVPrXrtGhy8
vUKXwcYxnLjZNIRlbaDYSESWFCk7qEpYUfSyspxwhPkmcKcdUEDxXq8nJnUqRTw4fWo87GE8M0Sk
lSt2BpiaOU3II77J/9O/7gMH3hWc9TajZY7cgODea2ogO6+YgKQOLieEg1FRQ8KdykPbS0MWsDXb
rDpH/0w2VorRqJIpUubGUz1nVu4fspN5BBJzDkh+60d97DsD4kz48MhLW7ozcQUKG9gl/utappvZ
YNMZ7dqlMSrB6ZA6zy+nQnxqyLojD9dp1mIYDb2hW+KdolkKMzEQSbJXJEb+FG+rp8z2lg9OTgjZ
KGTdTcA/g9oz09LEPesa6DLTRhuZLpGwvb/msR2DXSpaMeBp3ParWF1isn9R9hf6H0qRvpgWkd2i
h2QljcMeS++6h4cPsuTt6PmFsENTMhzFO/q/oCaxWLXWkNwVYEsuvJD0mR03U9mcZ+nZS0IoX+C2
jf2FQQn8qFz8TxmhccUoDqtBiYWxLARUexkRY0mKeJa6SjVhTsc5WD0GlLscRq6RFixC5U5bYFGa
+20pAgrZzPIno6ASLoZRGPzLx5Us3M35V5oLVtiVza/sDe5sKzIUBS4iqgynrRlhwAolvAngESMg
rylZPoiGHbFJTmpvf3pgvVorTnY66mgpc04aKqJEXMVl/EAX11K8gvT9HUvjGjB8VJ1hTAgrhF0/
Vcu2mbKyxYESueF5EiNcAdJ5Rkk9F8MPReAQYpCefeE4xYP9XSHk+cGDz/gfk4i8QKVR4bJoBZoq
d/AkyDksKg19pWF4QBM/FH6eleU40++P3PIlebScmfTXr9Y4xBRXgdbyChXhfVwcW6g6VZ68L7DO
9607aP06qRCgiDTuPNpNl/daKRaTjPUGb5Lm9FEGR+C8s6xaGmZPl9YHy0Lf0SWjlaV6wLnEvG3i
qmhTKuMkOwS3mOLsyvtxqIDa8YE82E3+DTvY7Yp2WZM6xuRY8RRo65rrdzpGQHe2z3UvPP6I2oM+
Hl1zAebr8LWSRhO+FU4L0nIAP7IkHZfBfTkV9ViGpZdG2if0EnmlyPx2QK07t9wFu5ML7dqLPgzd
DzjQe6KQ7XE0/HRoN+p+IHA2+252RZ3cQIeTCs5EbOVQ8BeEAVzcPjWmOYaukG/F8DINe6ALl19Y
wVbDe59UeyK9AvQv4pnye8GNqOxzjfShNoRXiFAb+dP/8GZeB643OYr5ijuFoCWs0X7X8S/zd2l/
LYN+o4auFgu9rSVeCI5hfX2QzW0L6gxcLOejjlXJbIyVbZOBMImln7KToCcxBQq1TG4BBIysbMIB
sHJfovYerjLfH74o5SLACcmhl8vI1ybpnqSy723Qx4z0yukasu/5PJAutZCrrqikVxyADgJAoBGC
wRMtV/9HjeKEYWy38UkDpgtsIgYBlDmr7Gh3Icr2OlKW7OetDAO+bKFW66Wc8IxuFGHcs5jFTZu7
/viRk1OlVZq37WqZ5dWQHRIttYSmRJ8tj5pFINARq0/gqA0BhFbzS2EHtVBSBCTlvXRgtD7YmX/Z
uZzQ/DJDPVDd92i1ObQdzpFD1XW8eZn/AVwIXu2W9FZ2UeF+xfVu3Mm4cYkuv/oNAeMfzEzPMzdW
Di6IwCfVgS/8kyew/ko8QWlW9j0mmsrMBIWk3gGSjYLB6vHr8k6zcJOk3TMNyScnzPpxemDRMdbb
xrTOZBVC444HKaTvjaWBSvTNQ+uRUv8QLyGqhHmiFWyjFRPQoRi24gCe6Nm/KBWXjSANyy1p9ZCM
aR0h2QTgCvn8p61+K06PEwL/szTm6hTfouJGAcG1CEaM6n8qbboFzg6yPvaO06pHatehD5jmtkli
9DbLsm7ig6g5ikOGzC1rhA2peev7CD0/Iu23AwuT8lNvjEVWzXAVo8MaoGTiuQacW0otjTW82+3s
fvuakJf2+LlhpYVRxHMV0dUDDabBMHsu59PQ+ZjlbuHBu8lN0kAhdnmHhQkdlplSPXS3QskrFl7e
gM/5EJd7wHAUGvQBcWtU1lmBBoF99alHXXSc0IRGZITd5Myz86ZeuDfjojq+KrDgv10TcK1A36/r
jMUxF/zAaUOLTBdAai1vnlqlWO/8Z2N35T+vJWbFuP7zWC9feJDX1gUShH+OGm540zRPhfHhyk2H
EzTdkDDLXfcte5eGa/Lh2f8ozCql35Dp9FoM/HLycCmYDhgl1Yf1suy/cZ5CHj5qnPQgMwqKQJ3a
Ex+chkNgtcsL6u1tMyW4S2IbXE+P8OoGlXHF1IDAtVRtmr4RfFeyR5ErKRldvN6n07atpQ6Kc1Eq
r1wfRoECaI14EMNa8xSnPa4cJRrfpHSWgr0pDv3xwI8zntrLrQfDw0nTfEtXY1za9WMFqTH2YUi1
vhu6KmGPL5xUxFUT+UoKJmG7x3+tOLJ0Qc0LrwBiPQEWyOwA9xXYkA8/U/xTd2kZ+ZM6YovUNsy4
7wPq0AFbQ2bUbQP6NCkZbP8vxGUoLMXt/VPhcM2DagPa352VJI29UFsOFd0f6uFww0iqpHDSHSWq
uzTVgXbRi7T/ZSSKbpKBrZW/Wfzz2AUhjL6OUd55Iz5e2FAxo2JCNeWm0ZDx6scWBZwyajB+mHin
miYjlUOrlzlnyaFn5KAZvMQDxWxknjHImRqlQEjdMSjn9hJuyDVX7D6ljGRTkMzUbJq8b3zUVbMv
FwNddhs+0tDbvr8SF96rOI6GXixj4ifsZH85167mET+XyTqXTiIXLweRI0qA8ar4CagO9eGZH180
6+YI2tgU1Kf9tO7Xcq/c/JYccyswF2vRx1//eElezRR8BjJhhUw2YhI/la/a63S1YFvkdAQmuFwY
kMGIDlCgYGbvo9f9CHVJKxpUu0Uc/9OHqNS42v5gPyXrSMmDA2TJFDQcIkgWYhITx2fIgRbOgEyX
yLHIo3zI3IuRUim89p4nAoTo/bUxD9iSouwsTlVvowmk12MlGhML51alyprfxTmF0VvxNFsOotmc
T/BKqtcAKc4H8p3dyj2D1tejlzfQCDwoi6SUA5pY9g+o7mk3+Nx/oWpEvWVZQbh5groQ9OGiv1DE
CG9low7Vk5+pZ7MTbjW+QuhhidgXnnSSHnarCq1OEH8SwYhivLxDinjW70SuITXUFjj2+apgiA1d
3QH3LApP6zh7Q41V2hQRue3/Kj0KBb64z8WKHZiHn44eXSx2vQSbHfey54tXI+rvG0QRTFgRP05H
q/6A3slA1WsJR27zqrMsQ4mDVuh+yTxPhVZXp108suaYN87+RFqa2YF9SAxkeKoUVZioQPAkp/DX
t/0j+DYXOt7khKv+dRdzhVskEsNosAJNGiem2rp/3XCKOz8fsVW5xTAVDXoEXtHneFX8oXNLymRC
maGVsFp91GuIlCM6jcwtDG9AH7kx3fQ03cHGM/tVX+tekOM/aGGPfX52D80VJbvX8lm3ZH0w3MPB
5QJ74YEEkQv8OM7H6sMIeFdayMn7tSck5WDeYNN2gmpNB+sYzoBuJGvgmoiZmQ+VyeX1qA48ysfi
LuFv5JmKDBY6EMJCKX3NCshfMuxvroQ4KeM/TRUcNR4nY7rfw+s6g4PFoxJISbWw2txY2PkpaB2I
8U8wWEriuKZ1A6MRoksPTIJ0sYKo/h0X359vr2uWyw03pPYtX0PKNX1c9WzjqB+zcQhfJPW7t5zY
wcHhX2U/Sw6IGdE3ErQbVYusxk5zWGq/rH8sc4QvHip8YSA9TTfmQ4wuYG4hauvQViRFq4aZE8os
v+09r85PSkS5I7d5+uRyIctNgyXCOgwZBme3+QQqt2v8LJiAcCXkjQwVShNYrZRF0yH4A8BQMY+U
1C8UJ6mMeYtwPMzTiuBRd9cONwJ3cTpihGWgDXX7gcjCCzxJVUgY6wB7wsrn94exEBOc+BFEydMx
bhWAwfrzseG4pjDSjV6xp+lgSoeH10tp/XWGThT8qByQFGILDx17T3DsT4y+KKrcBOc/tdkHm78u
VLH65PCfDtp4P4tOZJSo2izD0jJ9bpfF19wdoJ7OhKTTeo5RoevmliTq8XOmyJZyTLvuSj7+bBeW
tf9B6ps0M1laXlmu6l9XCWrzJ9qpaqJJSPnSmCEFA7cjGEbHy7/CBaMUT04ObbDP95OutPzatgfo
m0EC39X3CTZnSojO5Kq4d6QkmUPvA/4augV/HKStz0DpbdCRWAbxm9mGpQyt03KWnp7Wu342+U28
UgTBH5LehCcUS5gJGs2LxjihsahO4oA6Cza7uhrN2cD+esKoRQzUX+YFGarxmZl/25Ope4ayukO+
/06oMT0mC9Ppanli+SnLvAz1je2Q4qYlGeHJLqRob4FqvIUmaQesuoTIDguQf23Y/OV5rALojvQA
auWBy/tD9/Ez1TMhUbmB1VrLoK4ppMHV0RfcnsJcbMxuQ8vlsztMeT4fPFPbgoIiALNaxnvoaFdT
kW4pwyq/C8QkyjQGvsO/38/ZrQgea8Omk/wedyBJ2XaxoJetb7UXEaGROURr6zTQ85sTbHwfDJVI
DhZpDMzhPMH1anjfu0gSslGNLC1hyh5ZZEHxnHnWcE3IQpaq1zUYu2p7ltpHHF2ELlGsOMDLXWv4
kE0FZBfVJ3u54PD3L9nyUvdi6AoOwrpyhvT1tZ4q9duHGcPzxwPOSdP3+5fzqYNQIM7XAJZ5aUwL
55Uz+A7fwXk6A7v2LZmEAH+eO1LjcI1hLqscByygLcqsoTWCM5VFPlPlSMLPhdW2up56cO1Ldxfi
lqscqaUzqVZGBAmMLvQ4GoLnfqa0jbMTHfMO4XouMWRVc3nbBu9lkp5kWdVDEQrdS2tZXObhoif/
vWv67YrvHouWIPjTzmu1fPoPZpxLXInHlnXGJTpmwX/SPfvTtzKkPiVsT61RF0QMwOiPZTVAf8xB
IGbiHDYVW1dkg5zt5sNeUOaVC4fUA+ls/eNWlGof0JEQ79wPCQUcdttXF8wRVxH9u7xwRuM61+X6
w8iCTB8hENj5FtQl15wctJZ3zB+rUYVj6eZp7nY/wYA1+WWJJjAWJ6uCgIVAU5TCl03I0w9gVx7G
5XeUBqy3ux1QI7klPGRPerTY3OdyIELn6ssqnWGOa6m0qWr4gXQ0vJUkZpVLEV01kuD26ZHQbuOI
SkFpuo55Ge42VdcjwN56d6RY3YNmPNBoB5yus/a5EA2+GiNhRHg/s0g3wlx3IyFDMwMNgyhZDAQI
DhrgIlyOcJHjkhho/Kh0zDqiLJKVQ5c8r/uxNPU2481MZADYjjQpXfF+f15hYuztCG5I1+DSZC+K
pGtij+gpIWLOB+wOWos2pVtTNfIFlYyhkfIJD9hPLEE7AVTOl6029gtg2N+sLK4v4cMnrEymp27s
vHvSKQDdSUwsWQaWt4iALm7/TMG9ZBmYT+96+fsL7EwiAKDQMtHiqnDK+zEmKl+3zbf4XCFGb59P
SeONf3NaFW5skoQ+UsazkaaN/fucHnNOAVxdmzRHdM1UiCoy+HU/AC3qF6zFTdq9lzhJZm0dPlFk
cI2q7K7rP7NDI2qi4qQQmANgO2ZgSPi1WR+0077hp2YVNSGm0AX9wIr1EujAUI3y1I5S7PNHBmaa
kCDYolhEZgHu0RnBqL4GPhy9kiQDKreOjnbg0koPTyOB4GtjNZ93woj0FMF/E7CtHXjGe7+37aIi
aMTRPeCRbovHfWHozjbjbbsUOip54bIvFW+QOQZg/CGx6vuWRCfeX42YXSvtIq1nJYILSMUxWF+d
8Jw029J+DWcErEKz8kM5zwX473gBSxhA9pYWaIgCOvePWqv5ruZWNAIg/p0du6rufiFyqQmwSo2A
+mMMJb8HJhBZ80o3+pWP2m/ACaLct3AiDxrFQ9azPrnPUVENBTggAHq4ix99amNOuTgrlrVrt5l5
N9vwA69g0BpHaXFxz/0AgPh7sL4OUBiB8nHNCwpSjxZbpT6NZYBUE7xl/KZ5pLnZJd2mDlw4F4+I
Q9mCb4Fa2DQSmz7ciiGrDL9VMdsjexyrbN7usawvCaa7GUoAtwj9AttYYZeTq+S7poyeTIZPmi3L
kqdpst6KLeyTT+8xT4R3tvNDQH9UECAhH78xoHZ2D6F7dbtX3b7Xh6CpexruWFQ9SA6sYLEa8m/4
VTG4iiunMMw12bC3ldrL9/Fp1wKbbA3nVrOfCAqFChBwVajRhv5NjOjT5VfUDWZuD28cw4A3YZqS
OfXwnt1nJsGoMYJlI2PVCtVgISIjNbkFdGMZcigUhg1G+tsJMg1HX4GovEUKcvYPM4sJYxZuptJT
x+U51xPcXmzXCe2YctmHv1bl1t9z7s7T2B3UmfdHQvVRdU1RRb6cbU4RKXvVPabzQ9fPwCdL/XyL
iHfWn+drvuWJUhEotvjHvlPyPoLrP2JAR0j7s32fX4JQ9acqCcPnVXFNEcAniYfoZmLY15gdxocE
XzEV0Rsgijk2BcJHu1CP+H6ohvH9vsUiHT9hNP8wa03atgBsWoghMJlWEtQAZuYOfoDk30/M3+8f
EsILPjoJ5+ek47lwmVJjXo9RzxTk3seKZOEfZbGZdsodyivsJ/XG9nirQljDPppify8bipmchTsK
8HSsgEk6q3ljAOAAHQzrQQVGYJ+XMeAKV6ZgG30G5rArqhP5B5EAxKuQAN7/D/lNizhozO3DwId/
UzPvXBqVwQh+qni7ndbHvTzLK4LUgxYRbQJeJIU+N5snVU4qTaUhUvz9xD2aEviMT9HJY0qEeRRD
Ee+6AHkbmAosbaSB1crQG02Tiv5ZyBimsQBMapLGq+j5iJx+UuJTB+v7H/p+qzjjDXlScqB+PRCF
2br2GEP4EaUvCkZITLFXboDoXitGQq+R5z/dqR9l6WtDYczXWURuQHMUs4NHNtO6SSbgrqqiu5bN
YUMoljJEobQyOceLPvcdYPYJJkS2gXhSAFQmelLZncoAb/QQakigZUsOx1ku4UgyvxRPr23YryDc
A1YkDalSXtcELimT6DCcT/kCL9y7kzImwEDkPP/6MV153J3FDTuwdGikZAX7p2HyDp8oz0vWBsu4
NQL24DjCm5jA7eJGy3S4iD6vYkGQtyXMZ48gStSADVGvLZeWuOfnXNlicIJs/RKuBMdLzUofcHSM
8eAq/DC3RuYzJczoNRFNZDg3eusf9bl+QPauEvRRX1hKXzsBdpLAOdpBZBveWdmNRBJkN5yhQe0H
1XjSvt+AcMuoE2m/2h7AHn4WeWf1wfYX6HtRQ49IicQSht+r5rCTkWktdlUxJdrqGJEmtC9zWZd/
xuE0i8aRHw1Ty7xV0ZWwuT+PKVGA5kUcifxJtgMKIBDByriw/AL2nGMi+v7Sm2kN2ZRzhbJi/TeJ
K7pe/iJbvpnq72NyAlqh9lXk5+vd/8QAVMioI/agfZ0PNyWUVSnJyMh7T+lFJQ9CpRGHLrEblT8r
9lfim6Yh/L8nIv0zK836pzhhA85g6WiaQ6VBRbSWwYvPf22wnLBgUwhp+ak7hyxDxPGg2cdafNgd
njhsxw6XAMMzRMREstYu+BB9DmQfoD9cLokYSpv+XlSTAUxpz/DIJ2fIRccu5B3BvvTzEhwGB6AT
LZcuu6XVBnKG77vStVSPPFruLPv1wDjkYFtVesKlsYkUeb9rtChDR93+x+PKy0kZ/+yN0MIaxBSl
0sgCytet1X4eDdYxk7tYxBUu54MNmRhFiZju00prlVRGW2wKrpjVJ0JW6QUDBzdfpt/po8Q/vG9n
0SBMCO5At8+Ux+fuBkPqZosmDGtthjT7tVYxWSmWwqwR8G3WcACNXLHXO27CvjWwund1EMcj84Ea
oWz5Ou3YS3ncnHbg32dCUjmP1GMmPI9Vjxjw+ZT6I3Wy7wxf8/H5GQWyMHQNLx/9DR0We06fq0Xa
9tb90PYcrxCU0irV9v9p/lM6zsOV+qHg/9sjGBWt/+S764Vu49JbQhgjj3hrDKIuWwnVI+zi0nTH
Uq3v+uHeDTCUWG7yCoh8T4Sry/Itg2L6VzIGNoXjjYlvldHJ7NvBQ9hueWx4V325jDsDEh/pZ7a9
WHMHWZYPw4HxrLx/xpl/P97ECeVjbDrFAIBUKAVb9zXLdoBmtBgIJkw6lss3dakQFovnkho7vlEY
yEuG+Z6kLWO4WJGLBOqHni8uQccMSd0SqOu9LTvgDdtjT3enik7ii5VstWSIFfgVWeTRwqc6x2wg
/6VQaNDLhzJWmIcUqLztMl52gc5sG8bLsDzMPyeyMKTcel/OqeOfzEwEZUukzpiuzqyrbBLYyHCN
42JAXhS8fZU0DYdp33JyFfcazmudIRb23GPlqlwGa1SDoNUbWeJzwnXCeYYAZblJM+NWW+hUpEEq
jteo7eU2Zi6Ic8HvI3LtQ84lT6vl5eOIx3n2qh7I9p+WIqeKjNxIUyi7/x6XwdoR+voFDOfjdnPA
MtnSLPTKQYaDHeKCUSF3zI5rEKM+mLCC0SOz2JGpvrC49ZBcFlcNwSj6JC7G56NIJkD2eA6XLLuG
RUSgoVyT7C76YzLN7jL1oxb9v7tHGVZmim9/B9K830Zj5SQi3lN63El55XOtz/8mbvG4tQvydnI+
zoIKpAH7FZ1Mg2ljxASGKDUrdpuioBpHY7+tHgYNu6vvV3VHpAHgKFrk8CPmc3XdRdwuE/s1Q0XI
WX4Z5IQMQkOVKYrtJgW87gkPBDQWjAzniS/P7K+d0lsanXqtZ52jqBkCw4oh9UTdHOWph5DYreli
zzDAehvEGhorIaAN4bz5dyX0iuVsju0AytTQ090YNNF7YeGPz/v+7wrgaYkzu9F22c9wtxtR9lTx
bPZTh29hYA6hLKWITLXQyeNn3uQqB2Rstbz8ccZw/YglqK9jYqh9Qf40tYv9ON1ze2V7LNhSIuJU
2k53P/OPZQ/XC1iYCqSewykFLi7cXzJRj+AXF1lD6RqKB7nQdukpvNYZz2dosis+QiwyGEOHXEIR
8Cgc/5kanqzpRujrSs9BKDTaaeV9yNVlVk+NDTh+1lZJrPRjQ/monDg0jaGtLa15uzmZe7ZK4tbd
+kFZQdnL2VqGM/4cIXyJS3mU0YDPE0Ir6RZ8MQtbdut5ZPAI81DpN5hgsnppoAnP/lpl37Guc98v
H2ZPCTiqlaUfbjHqnXIoHAiDau+aYIOB3yfLAf6GLQG2eerPBAs5C5h955xZhgb8Hsfl78GdTLWS
NhoCRTtNobgAwRhllHHW8K47em6NflElvO4jjmb81xR0jbLOrjf4gmBWXoeBbEj5rYpDLI3cFzXx
H87E7MdAVM9+mc5wx7FXn0dVv+FjZiQw65ZLTSVc/2B3qgOc1QbrCrSJzksTHu9FehlTjORcQLo/
e0vVDZbNzopv2KNjbhBJF3Qz5QzLyGkliBOFOmjTnWFnKOO7JcmnvuMg9Nl0VYbfF2pTG3LO5VVA
6mQeQJhuTI0Rg7LnKtwNBXY7obDQ19JLt4epWjq/tAr8HrYyONbTYBqxfpLjy40dO/9EEmmLSQs+
w2jSZJJIvpYz0MNYJCs5qSEf5uiYcK/wstPz/andN2pGXz/6OS8l17cy1AgBWfyuIRYORSHkUE0w
Zl7d2s8zKCvkctzSBxsEa2mXX0PS4YjSU0AaJr9s2E1fISFj/ZM/MFVWwjrixi0a4wjC7i2z5Dib
NB4XkciGNZq1w8NaD2vLJwJ7sgRBRyL1w1Bww1bE+nPr2liaA6mLbQ+IRLX/MVu8y7mXxG/xKHRh
eeXZY/62x36iP83koDiaeZMZT9xLv76kUAVxNcv3/mTSf0TM8R3gyPegG08pF2FZouQhZf6Oel+s
sUakznwc91utfwGZFkvIiX+GYOBp9BT/in/Oux5AGhx8GIdGl1bn3r5fkM6JG2dYLiV/8W6qHKDV
8+QZ1mMJi3Tpam18/MQssnF/Tjaueah9LuMHEQcNfoVaL3u3IAA+DAgbGhGQuCYgVqy4XUV9Bbsb
GEXDQpr+iuQDJSOXucTED2xBcO1mXgrnHySIABuk10OJIH54F05qq4AFbmg7WWfpnXsJyKhCmHKs
6eamjcYw/3TEBFOxrmXbtv2h0DhtptOhNS8yK7k8cD+TuB7/31QEjJ0h2AGGqG0hf7LBsiwzl9lK
RqDVxsAVgTv6Dl2Glyyl7PR1Rd2UNRmLLdUkZu8I1nxd6hOm+xaO++0LYu2lfLqWaGh4zfCGJvsy
ILlIcq0a6pawjZQPbB+KNL92MsoWFY/CA55iU7TSCWOeUK3m/QCAlZWVIcZHwYoEGA7/hZHX9S/s
Vk7D1eKgGwpqps8S0U6nlepGEv/ku58fYOIzinMaLZA9Z61pn95Lu5zUUKUERqqIUBUVspiB9Dhu
KkmzeXAuD1Eqgt7U41K8/cvwZrF60obbShsOPW35JageMhyVLF7VWEJNVZb+/ejr8+IPDO5yOQOO
3aPPYTvrxOKN0nHZP3ZhNGkjJbUUax3ucSQB+VtuhY1HLC5fwPkUFQLCsmgC8iqZLLz4KJyoPAXw
iNR/vZELbfDEjP/8ijN7p5iHS6GKMA3Ss4TH3C/wP3QdK+UHcaraeEC91juAof6f/Ch6T4pGUG7a
KULAyrTGLagQFy0peDYUBjnAmxRrNqWZkhWy5EF1b+kNQFRpH1O0Uu7ofTk+WrAQZGSE0j8DRKRY
fHMAELfdvHUKytSHLg1oyADu7ypltvm5U0gi8sloQi9W8JqPgQevCZ05buY8j6kc8D4Cjn5+nBLH
LhcyAp/L91x8JdOp8XGwTrjQN2RaRvHWozdQVbIe0phEuPNoMa64IHHkOLVqLdpfQy0m3P4eVuul
658xSCSXvirFfcGdp9B2eW9ohSen/voc3Aj5GLXRa4U634iGBQIf7PMaUEv6KNtxCW5iMr4mQnaF
jn+GrNhw2e4a9DAkSvYJ28ThLYo43KyAGwrn1ezvNLfl0q9bTP42xkoXVcV/602fcgDcCn+EqsVO
c0gxkQR4QKyxSiXqnVD2qyj9lLLSkovQywHa7yUfYWDwhuIZncRqdgNN/8po4COTLs/C5BAyzlgW
f14LlSyqoWJXWjb4mA0k8cm8oV7z5y1JZ2zRuurKohhAT8oRdso4VGa7J/Uwzsf703CQSi0CEY/v
v57SMyuLlN6zlnlXyaYVubc33nzKqfAHqQoPUUnwKOq2iN4XW9y3JHtf0S0DqBMrIg0PEKpG8nNy
FNltgvQ0XCc0BPKcoFbppsYEQroFwvEbykEU46T0gFKxRQ1clAPIIolwKjunjDsjyXmqOty4WwNk
dR+ChbSfYfC2qoJosalWpJjJbCksnlVNgWvqICAhK7zHp9qPnfk8coT4tXqHdmwmfr8yrXG0Ezpc
mkSBUwowurh/8u5TKQqKJcBruDD/vOrbvl87pvlTRH2S0oDrGSJRvjGSSqwc1V789dQzjP3aUPjT
2VUAMOeB4tuaNiEIzGfqR05oz5cBcSDRBNCDTz4JRNUSypIoubZIwrT+DQ7FgIwNnK4RALaLyxDq
tdOYMeMA2GfRKSyRyJ3qvConmnEbXXRyPgj/FxUVJXALwzafYiI+fZ0rCr1cSI6/ppAmrdeHnGfn
u3+fP9vjWeC+DmjpZvFApNPf0V5LXrdk0PLHydC+cxpDRiTOvvFNCNYkiyg6pClYfnwxk0eg8es6
dpSAVV5Dmo8RzioVAKP7G1VHDYvMlE85GG0N2kJAtu+O+ShkQzCNh60eQY7yuJMhp1thCGIVzAAB
y4VC6983M1QO3nyXNC9sd4yUNofgfY+n7NVjNjwkBE5w/CqjI61QG3A6q9U1tXUYHC1lxjYkUn87
rz9FJjXdHU6qhdyoat/McwY8hGvBrpsnXPRIB+AnzQMO3Na46xnwS8cM5CDquI+qQ1Q1ew1X67oQ
rXO96p92HZbCwMCIviXyZ7t2H2mC6dpe599QAsQ2jEkEQXjlm87KjQivHQct6udDIkvYX0kVmyLJ
8r5BLIE9WfGQr2hl2tVsCiZ7TcD0wl7UODa78y3wLiXzx0SWzCX7epAOFkK3iJ2d2UYe3w3tAlpJ
t1qKpfCHoabgcc5DH3sZUgYbmUMBizRMtebr6jbfu0j7gZljo1RNGfn9K6nCpd0CCPPvpPlABOw/
eCYwWOsbZjSGUUtVIXO8Ux7rj2AA/FlP0fKQtbYpN4TOGQzopBHVtav1oK/Oy7AhYsWKkxYIjks1
gnkK+Ok/L19iIYaHzWK6cCp/mix+DPof+1LLLgy8pHFYhxNLez221S0LfPp9GeU8xdTweMhSevsS
okJ4TVfqaMtg19i4lDFD0vgJSpui4Vza69i0lSiL1F3wLT5lW5AuFJxwc2bEGt/iFAXI2rX/sgyo
kR0TaCXM3dLkWBvLJaOlm1+jirPzVDh3R8XfMNzfEmrpY9VZIqYU55C3Wr2Q54vYUKrLp0nXQ2w2
KMsM10oW23O5xWuC8kkva5QZ0br+/yvas51IMG8kYXVvvWRpd7GuXb+e19YMHipnIgILghut3WUt
gDyaEW9WCLMe093XvGA6xeBj1w9mXkJOUjka3chE55LBL8nA4Ihtesq6GpyhXpFzFXeY6GuK/l7Y
8gpigQAsEzj6P8vAlAkUMxmto7ep+ChbSoJrBHEGr28jZSkEFIkffS6AYtl2fccIKNczvkLcHklf
VdvaeZ8ToQ/LW6ae/k9Lw9QQq2TxNSHW9K1dZpTURy8ERFTZPOEg1FUf8dbW6YKnSZxY2GakHVEu
tCmvjwcK+oX05jMwszW9TVaNXS9hKcT9hHrDuqBzp9IU4MxftJCNE6Old4WIa+MDGmSAYK3vxKkS
I01Z8czfS/vF2cnljeTH879AV90C9BnyoDJqZxwTV7IgUgWmYZRCztjouaSZgIBolvo5H+e4btfL
X6897FT/z7yRjNkfOYOb4EUPseeB5xg9S8Vn+mBJBAyu10I3h2nz+brJestPPL9+lvZ0bIV2YXqR
hNjRxxGuY4ReCgY3PylYMhisMXcX0h62nTqPgi2TEBYFfJ33IpZwL8jHt7e3gGXejER2+BGkg8OG
fMAYyMp8pAiccydbA44Hs/Vr8zuMxJ3fY/LyEXgF40EwPzCRDcfBh7LENQ2fT4XGoD8jFjmvVDeh
8nWIpT6EdYgusvSUK+DkYDu+1XfYMllGskHZ0/VGqGToXGnRsGmMpOqtLyHuOxoAG3lqZhRFrNUO
w2snRzV8O/Gr1oi/Sj3laO8BNo8xp3VsQNvuhAViZpsQevNPzrQiD5rTryYs2dN7idiH5BMly9qk
QCVgxzxjXlcRzNfJyNgOxQsl0wso6G8K1EOyzmXiMiLEooHnFjrOa7LaUJhjFKhoVVDWh4BvZIbj
gLXhKKiuvkqzufiptvwurcGb3xR1lmRHuhCufKVym13lde+WTXjB/7ocqw1n0UDsxdOtVODhxgjp
flXNW/Di+a+LctOzOeEXyO/hHIU3vkdv0wQfhkbsqyG2swQh1q/OAVCIPhRjy5K/c6zMkkXUcdZW
l/dCWUwrmkK7K41bYXZhPOzn8wPMKPXwdZJcX6kLc8P5St2faq6D6la6H0yyRrvkC4CoKK/DL9h4
rzZTkUQQQzE4UHoBPjwC8HM86kIS/QkN5OPGV/TN4csxZazM3ncKt6/CCcWZLZFdtvBQMAYljlSw
urBqsw+lKpWWL+/sCNnkIXLKh39kmQG817VI0IVVrnSvvGJH1b4AJxDxbK7JMivW3aeDSlwOwgTH
ABz6uXlFlf9McVEsZ2GRN6DXbTJikDViezfobi30Mjhlb7MyxZiYFs5pKJAs3szJubCDloiMG8nv
ldusvKmA2gcTlnvVGVyMQ4kny+RGDD3oTXLuIt39lzShkyB+JUm31Dd+bTGMA4AqFcgvp5bBRU1N
DZSM7a3b6B0JuPxRd9qcvdSiW5AYFHxWoi/mQfvmhzJt0VTyXDjLN48jcK7RmIX94h/kxwL4YyBz
2LSxvPNE5kWAO66x9e4/7agqpkNVpJlMSlojYc0hrMO6v4FaY9rB/kPOZFWHdmOCiAl0U9gTk17o
NUF7aGwKynX7yb/44rzVEh6F1gJBMuVRffpLzVfz2DCs3xNR0yJgyG/f8dXVtBmdDZ0w5aaHeAsq
Mf9/WU7rSSSDG10JLa7udRj6Mvzkv0MzEmIX/L1CEBw3nnbPOQTzR8E0fSr/0AEiYOF8z+Z0XDVy
Ai78xYxmA3mwGGnK+I3+cAH++/wyoth+hTGH86xVFeYtohbFDryve0HRk1Vl3yiS7JvdvLfSWSox
x/sGYcDLuE+tT/tyrC9n4zSoJ7RiJBFOQcCKLFofsEcNVOlV4ARb05Li2UNBr/H+jwBKYDEqvx47
cmOMN9Y43WH1+F/mU0usQTwzjj5ZNecUORflXcwwQaz74ri74Ic+8CYRjrmwUSJGJCS7jy2kgOQ5
+KfxIKtAera7gsEy3dnMvr4p3aJzHewjIt4/GPKvyMfXvRw3wRWHpIay0RllZLCZaQ4zp8RdgBR7
xKGADmnKwXbQPNUlV6XiQLodFtpe8rptnPehFe6LONOj10W0xAq5ai9aSXjky3QYTsO/LFn0OzM8
i3F6I8kzTzF3kYjUidXiGjhEBfcTJ5Du2D3Jpi7LABJa6njaS40seLoLCDKoLdGsgv42r+2KgZCW
tyLDPWwLl2XzM1wD6bEdsnEGin9/CjCwpnEasJ80Rmjw6UE59XB0cF7BGnJ48bnZb8i/vqaw6KGU
WmbxZvpEehWgzm2KQ/E/HKFHHz7byJ+pwT+8cK4ouwjxvZBxze0M4hSRWlfuKm2iNaaMvsKG2kN0
dr+VK2+fEgvI6tsciNxdpl7b6KHZJDMPGAra9gx+5zcNLheVFH9CTgeRhzYPBdNY27uydsBKuBWZ
BJ5clJg7xpt3d6vRYvEpAzLHqY4HJlhAY2kzfs+xpFLvIM2PbTY02lExO1aV6QgSXhXfqXkD4Kd2
dhw/5r1K/kjw6UuYLhxHmG6oBNxM4tn0IIRPK/Gih68JCod0ghYxyeGvnXewVx/FbwnhZ5kZzIuU
pTw5bni4QnLJwGNdnXSbVwASURx5i1UpVc/KoM91ALVmVD8d9EF+yCz8NhL/ScVeXy2nehGfawKY
HnB5C57Y//7pQEaQIdBJRCqOjNQ6F8s8YeP3mD7duHy03hX4x/ur+6d4yRN3cdeRRRsat4/OVjJi
LN7c+bXXoDpHPTXkavsmphYeeefnyZ3qcwiAiWvfgViy+pabxCZ+YAahj+P3hqByKCDLyZNO0Zt4
8rSmXmothODF17eOLsNjbGfO58bUwBCTJ5JU98AlzIZdAYRohewakJurMr7zVBwEMlvL86goTbpa
DxMuxPOfrL6MVQc1FqmII26Djzp5IH8mk/zQFKniYNtZLYHLLPANsarnTGSsLz/nxndik8u2uiia
9APsBD7KalxwtaXkqmWtMghF1tLUdwtf7JSDz/hOY9p+xxuPT0J3HbLJoVUMrI2sCM8vKwamaoKl
qJyKNJfYnTfheTbCI0vt+fqFaztKLaqsZlIlTxkm4ceD0GyZAs/SF688OtLERta+6BJ3eFPAlkdK
QdSSTW1HziujswqPR3D6vC+01ptH5xGX563MwWQDtOEQiWy1bMvlQIka5T5LRE+tAKggSro0SQ0C
u+g6m3GbjOZD3pMRLfmXoQKCPSho0lzHtaV/pNrwMNonYqdN/vkNtqPLp/7xqNBcu8k8kJNdjAmt
YAhERUy3tTu0rwIoizvDc9QjMKutmqKU2Vj2bohmNihVg6e3xQ6PWbWGG8uUUhnS3pAC6+bIWOkT
vd4boqQUkSjMVmwJAWDIds5TpIYTvcIiWLaTBkikmd6FfAU8HZhp/FF8c//cKag+0x7n4dfgbE3U
GfKi1ABp5NxeMlspIlT+ynPrgcS6QYmagTFEYvBPxrZIL6Rdezi+q+qi75wGc0C2cX30QLxnt7ca
hoIfLCWjuUcCyDTVIVLiuQ6yi/oFkaWUNThzUzqZcOjj6mNvXjksdYe1EQ74OHy3WoVeHHymjPJ8
7pBO6DoZnvWy6riObzmyFrqyipdf1eL8KHZaKw9eUinqodiPGCoUFI2wvNSAIoD6Tuo9NwMsoSmv
uzlx9uUZ6lQ6omM9QgrahxkaocAEyuLNtYYT3v1uypOySd4xtQBj7OjtKItwonJuTIRqUPPbhOVY
outowN/uPmE8RcuM2ErHKiW244IwCKp6yOpCnym23UOVggIl8xmuHSxHTUP9224XJ8v/VioYSX9t
4kAIimdFUG3pfJL66Jx3EwTOonJZqL1SnSOGXTBibPIu66z+ty+6VJCtmJAY5uR5ntzUZdaBpGY2
gDsWbh7dw1qohhW4P+gsrvuKl/2qGqZOPHduKekHJ2F9yLS96TIbgEbRK7Fcrr0fVAXkUw9ZPw6M
Kv5WcPTtkw7XxHXx9LEUkmGPVMu+XgU/5mgFriR8uJtrEn0CMbK8nXGoK4d2CgdEdxEsfDDHlyRS
Zg8G0al0NFIY9wBwAFoHebptLHHu3m3egDlV1t4Ia+X04aDoZDzgInoY4BQ96Xgo9A9O28uztDvR
7DmSudhvnzALXYQllJ7+CrCKC9Su0bShg6is7tzfID1aows5O9Tcb44G9el8TfJXrtYrlp/sSX6f
LCF9938j9Z1X9nJfdNsW0XtNthdYv6OJNDa9ALHBl9q2yikcLqUpEtW3W4OaeXQ93PoNrkbX+MMY
hNsUEy7Itvs429UkN8j9NhMw/ioheq0GocDELuHGqeHVcXO4sKwoon3ITf/2j5e1/yw63EcuI5YK
ijJblWMqVu37c/bQcCGal4A5FGgVY0G+9oYA6k2utjbOW6rerOQ0IDVCtuhGB/mZdAvew9DE2Y+r
IPlMZefvOn1hPFd7gS23Vr6/A3QiPnErgA7g2ASpGYSFhJe/dt+oNnB8tpqTVbzTdVjghCpWPY2E
8Bszj+EA51+k2hnX5MGAHFMZsGYeJeTresmKauXpRvTY2HmVJSKzXiMs3yIP5UVCrOto6EfeXKFW
HiGjZMn5bnkV5NIlfHuSeYVDG7Jhvwm74hoQWy1A0Mb4QbzgDM+4K2Ffx/IfbZCaDbNiY/zY6bf/
yqDUrF4sF4Cidme0Pj9+PkgKcjKk56k5000dQ+yjflgytaDqXJKMu9+fujRcttm0yUSg4Vdpc7tv
Jj4sfNlSh191QJhKST7FKxJwd17H1iL2nr/0kslGXBDT8w3lfsxfEEkz+pHchPUPWkoMoEAg1io3
9n6sYgdSIaPgLKWuLrdrijjnJ3CwzYHwCkQzwlFh1DWY7c7eqsw6qjjCmGHnGzYLfxqQDyCPhwBs
XGmOskSOO6J39KnYDxc4w08lE28+ysueHx/HaS06ZOMEqoWx57A7m0e/XTbD1fuC0gog2ytCKtHZ
nKE4DPGkuPIWEhrytQvWnmHhPt02oDgJLS6e+sw9RTR6NzGrj3SuOw75GJ4DH1urmI9ZLsqGgVWR
DW9Hy4hakVEROdPJ2nsbEDL88DrLM1hCwjeAYyV8cBqeR6j2C8LA4nHnaeJ+5Lk6D5Oyc7QKaCUL
aeXWVMg03xwIGOa6yQjtPZNO5oB/iCyv+NE6vhevSLWWHf7F4QilW7NPj9WAbMFrHyKAbZcdMPV2
GNSkpTBuXpLdPRKn0LFuL/JpYglE6JCHYndtaqieXtsJ729B6PN4jf/i/kiuq6PNw9hfIqJYtJQj
UMiXmBXaQEYpgQjtjH23K+pa6wYEN/uZXPoGEjUqdtvMD900+j5nfEpmGMLZgIkW0SSOcpF0yes9
lpR7frnf5iFdlyvNe+Rq9t6GrJg+baaegLauR9wkgwqj8i6mrJ6eomck4LeQgJMTlmMyqaTqg71X
BJ74PkUaHNxSOlTWdnhRYzE6Wm3VcAW6/0nwx+rZ3JuEtO6nEk+uYDJwu0cm440oLugigt7S3W4B
kmpYZNWtH7F98VDfmoktCIWLBbfmqnTaisxLrxKf0t9g5oXLtFnwGGAdyT8urM5LRGEFow/UPYFn
sF3cYiKViLfW22gvaFGOtuNZTnG88EtcPndKHOo7Ugt1H0Xq3F+wPf0oeIL4JZbUlWoHhY5Js8m3
NqXMdyNaTlUIUXoWawGxs4I1K0clWZtq1ws2U6+50bkYZkVUdxz9V7YDJiFVDryxaxTjeOUFFoPs
02961+4AzANhnXVbptTKmOhMViXuYP9wTEbHSuxxAGE7NKfuUlcr0s+Siij2O9qmNeuSqc2VzDkr
p4p3SwF9u8MkGMlrta/dj7x+OEHSEt9iRj+305HZHDy4e27T0eflMkGqCuKnYsvi26AneHLWGhOd
UwgdPGTbKGvC2qpnSAV7WQrcYzzD6IOo0h0A/Zq7cIbiT7R69GdTlu5owDHdfB8HZY8bWUwnj/Ig
bRaNNJvx3MNsOi80oAtJ6apHD66nCdVSmGRRQlAiBZcisZ2OSNV85/OTZYAV8h91V8XGQPScjft+
YJQNKqsakPNuX1k6Gz4mGM14mq0+Z9+H+MwbTF1xW5TzqrE4Tef3++e1b9/xcGG1MvJVdkcsJGSN
9GvT87zIlmHyPVOFIo6wuKvsYINdF0BLTkOBcupkVmgrACK/jQLr9Mz4/bhgvDsIEdKxXT20qLkC
+hr5AxH4iJrAeM9DSVmYrMVzHM+BqRg39x3LDRe3evP5DYeetPOsCgiTWS3pdaeTAnCWtb5o17Xh
cl3jJBxwtnqLwAtEyj9bszFQE348wuc5In8cScDt7oh4/K2kAPilYlnJC4rUB6bFOaytCNt4/khL
KZycb74Av3Lm01ZwfJvGNc0IX7shXb/EHHu5Uc0zRpHG4ukLG5LCeuNdrJBlgkcCYHmjleqTLdD1
a5AEHroAcHRlYJLuEeT+MxuXNPls2ADfQu0OQU9oWgsPzMLf5Vnn+KagWHni6EMf8ko7taF+/R0E
T3AmACaHuuy5SV4b7XwjS3YgIT5vtiamHCwBFhGHew/xmI2BE8k8H0HfR3oQvp4MdODQJXTR0g1M
Fhuy3e4/qMVpCWe3SzsEB34JdafhukY05lzFbxoZltP+zXFn6cTpyzdAXG5teh2gBZehzmPRC2xv
iEQYeyuwSmJX3dVwwF8IkohiVucvGQPQkt9qAjob5eOfKOep2bZnuSmzgJPqJTqMtH6KVEoUSjzD
Ls1ljKLprCJQ7OPfIl+XtklHv9bI/2D4o1BfRTmJdDaZKEsBmTbsipRBkvzsDt97Pf88IDdUHFP+
Sy2yvd7bLywjJh+3RfZiMM3593VbNUstSLQqaA8cHV5WpAje0g7vBoT9cfrskSijj4NlYC884uhh
3o/CI8KdjVUSjUJkoZHa03q7YWjrlYdlm3KYrmLJbUq2gd8KXmAcbzW85+Cb78L3BWhWS0MK7oms
NZLKlb6R7DKozB1Fk9/8/H69If5b7TSm3yeV+S+W0t5kM6IxbL9psUqQ8pZOX/lsU+z67ToBw3SA
FIHWGVIwFh6ByP03QNezPtmfXaadccvGbY4MIyjxwSoxqFreNV+hLuHW0abqabpAUZdeSR3fWYl8
wDdgvfRN+fONn7hm2XdaCGZUSkd94f6UundqIcpsoSNBe2G9smastoBm15SVprPLZUjNGf7Pz9li
p5lPxC5EScxgApEosDscG4lmcG+Bfb4slDDZQ9EYtNyi7KCupq3eE0NOaIfEdZmKxnaXKJ+Qg/kT
MGHpwfjWsaljl8Jrm+IGlf6xyDGlEIGq77ujvG1A3F5hwrweiAgzdzNB49BtKcKlOilShiDXbVvc
nJQDPKk91NZywWoDE/0pBZxNaozFEiK2UeKm6SFO1hZw0PReDNN4JkCANhZW9CzCU0qIuy5BMO5S
Jl5rNi75pUbqdvyaJdqqTzjikwt/J3FyKH8FJHF12Xoa4gsFcocucfneThTJ3wuC7y0UaBpc3uXQ
jlLu+gIE7ywsGQEAV9tEb/MRK7hFdsGiKnpGab3rtpa96LkRa2yC8azt03dQOV8oSp1nU+7eu7KS
JDsIc/89qKuWsgyBCJ+pXggLHYTKjkC52N8e8Eney7J1QLGcTWF5gnku0A1dnIjI9I525hlxPL/v
wHbCQfAakV1bZsBkG0psCLDCju/AKaBz5CgPt8J6X6tJfZmXXjBZ3bWPjf64c/jDSFbpBhiffkjz
lgJ6pEV8ivqj13nSM2iH0CGdP6lC/nD/wiXz3RYiK9x6tfEReTvLMkUbr3wRyFPuzmS1WJGICuOd
7dYINhTdW2ggjSeZoY9OZL6vFy/j65qZMma/M8lt0Ny56hzGAii8w0MN4zecokibwl3pz1Wu5oI9
myasiWfA0JDo2yBBodvubsF5RK7y1win3tNJDxMO9NkHGIXWXsPXdytqSQnP6vd8v1keZFyy+1f9
tluxJver3q4rOuw+X32aUMJcdrQc9QVwse4ibgvxukBuh4cPHSHR9uU0cjl3dAJfUHHYBbyG0yTp
f8B42rmegwiAEQIdb3XmK9hw9YCN5gMr+DejfFQKSBwkMW/SVdrXVSDQDLC3uvXKCnDepkc3/COf
l0sGFF2CPpussazjx7mOVnacBmM20tZ4+hfDty54frfe2gJVeOU0hDtIw7ca4rEpQ+5E5OqxoUD4
+JyUpgp7PfzspTa7lvDCmGiQTMswqpmWieDPuxfvPDL8evzS1wswZZsK9RI2FYi//9/RwGMyj47x
f/xq7dnuu6lTR/dkkjec9ZxUiB41fI1J7cmjkRXcPk03s5s5yeETJfZSX+IEQuH3FteUDai32b7F
2nBUucPnxBlqA2BTenMw/+gTNlxrTGKaG04fUOCcgdQ4baGvgeuk25VBHbYYxt245xGpLFTphNnY
9LLg3azsAItcETBE6NwlDPKrjXVULPowGYw+wg9vr0uOe9MLbQr4jOwAhTJbKZI8+4AvlgCQA5Bm
FLxdnEqXU7nwEhjlVexzvHcP7t34uwyJLDiz1MsEvJ+RUC3W8kQd0rh8y/6+YSO939h/6mqIzdQK
rs9TXN0VjTN8NO6cQkYUsR0uywat7xcwQR2eZEh+PrGlw6FtCvixE2y9i5xGBfgc3CgcwNjcn6GW
bwVoxh2PiLUOC8XUO6LBKrTqGKbNzpu6ZS2LsfD+l188wHgqVgWtRlPzYZBUY1KLvwQVC1j/g6jU
UJMnLmBJJucWmjnYUZkR229YN3E09i0fearuUjvc6znCnRM1iJSnLkab7PONJ4Y9mvcKeQ406wNb
0B2kVs/v7XT2QUN8wH4iLF77CUQfrydKoSGMCAxvfkXl5X00Itx5TAYnMWponwERnfsJN9SijWDM
xRCHFKhOWxR11mOvRRWbCjMKVl7ahYHF+92myaOg6+V+cEoPslCo4wqhnDC9E/IrVYhnZhtQn2yI
E4j9my0fjvptOBcC1pwYZ120Yh/rpcKR0qsKPH7UtuLVaKACAkY6y2Yji9vRPgLe/DClz+vtgobW
R6DJzBtUKuCdFR9cDVx8Vm98YmdJVXbpHVloLFQ7NPsj6tqxf0gWl8IVWo/wpfmxLQ8cwruxBWdH
XWk5sXPF4jR38/9205pUZeacLYAtkLZGP1xiemIbTd7Xh4uWO3rBjB5h2SBKwFyBaXQEe7fz8MVT
fqbGl/gaB4NeXtqM6p2h4pPIiW+v+uWWaAhhQ1GNygJtw5efJC0kSCRptNIpYrkB/gKo0IRuaFkW
aG09gkDl2auGhR+cjTirzhAEkKKGJq6stjrECHbfnb+QLGUXC5ZtiNUCxQ4F6Cp86LTWoUSPJNKm
T3sGnPNWRleukBX8gPac448d9FyOwCvjeNH6zakeygOwFJHsdfIkV4Yu2HNy6SnfbInucWfWj8SQ
ErmONgbubm7vhFTm5Zke1MbLea/7+dfTwgGCQZOKfkmauW7zgNkXPtEV1wglxEFoIH9vs8zGWGhz
x1Ln4erfu6r8fYBtOKB2w8cSdoQLxeDw0uqpe0C2obuonR2N81QgBhzsTpeb5shrTI6pVz+DAxyO
BXsxM+MLMs0+0B98Nfyw4l7WT5L6jcRXCDGWb282Hk3+mmCCbCqgviLJbnCwhF5BFanHRn7ZgggP
mTMz/f6hqoppHrBWPwWAY66J2AymGQlQRTGTrG0HyjVX66daWFVQwZQKwNq+QBc8GlSZ9K2Sop9S
C5PZi3MiNjhu8/AXEokAClWuHwWnTAgs+IsJ2paYmD4oiQ5l7bi0B16PfZsa+MDlDr08VFSRzUdV
PDwo2blM7EbpsPvR5hXJc/1pyDHGUitdrETWG1Ffj1Suh58bV6qiKjQ6vwFPft9J5x5zh5WtA5GE
7N2Bhw6Z5teywYZrUgwsYKl2ukhQq+SX//iMrfO5LGrj5L+IXhorjB+BAGUMC3PJmLqKcQPl7LV6
LGfaecqF0tvpQQ2Id3bGrIriannBXw3rMdQlkFoVcLlJi1zDq9Sr/N+KfHHQspPIp4dt6SiOlIgc
Sh6M59C/eSXSh3Hc6fuw3tCOx9UzKegdlwj3NqMWEBDDsEVp8SwcqtCPHdTmpCYynatjRn5JsYbK
w/KJ/7zGq2oYVGY+01B7OSbVro4K8jzSAPjLoyywnYkn9/e5QjjhnYJn5fBQvqTrKDSt4IyQXziy
Mp/AEAVhhI7GKTWOp7nJXUk3q7HTR1o2r5IFH8gCNJvU1pB3EDpFyIJCkpn/uMjW8Zx3JrA9Wi/E
VruD3IIF0canSmqSp8Mqp5IJblI2IRJBNQFBLEvI3EcaLm0X4KJWznlKwka0A6m9yke5yy0uETWF
4BMXh2ZP/Mqyc8rGpM0CQk06T0de1x0rENQchQ74vOofIkwSj9pe4zaot18sXoT7r3JBNSghq6gz
M89oqUGvar8KRYyJ+pdr3uCDaEw++dzyeqtuibWP5jTM9n+Q+n9OxRv7kbFA6c5mwl+ya34hmNE5
1mD2SDnMJL2iAVClDN3VyD67cYnq3qoGnxLMApJvq58/kYZkAsOwOtsKlR6v7P6bLqZIDmDzQ6uS
+Q4Tw3kcNtzEoAl1i/h3xnLWcLGWFvQjFY/7jTkBQNXlmhYEaKvE1vXa/5JiD5EqyLOEObvAFo3w
odPXznaM2usW9du1gmbQljNc5EXeT8aFYLP4e6nRsg6sEa6GE0Rrh606AgSYDX09uw8cENmLSh5n
0npjORXoW+54B9NWWpaZr6aTmyCJBjEEluy3Jvac/Sj2O+GeqvTtbweSeEUguxHOBBUl7D3krhzO
jwk2ZzQ+AQ37ArnUnLdIM9Wzh7VzWgrBCG2rM+R3/SpaJXNgBKrTMiTdGQ/VvdSjH5xDypsGiNH/
Zij868V5qQKaErt1tl5lj/ZMqvYBv+qZWwySoXJJtXDDZwMgPJxcBD6CVWHL7xxlVcF52e9v6LH1
ChPdbDmY/wvMAtkLvHpOSbZ38w2Dlns4Mlv9opM5Tc56d3pLW94wSufQkfncb9x5fMj+Jh1XRSYl
mvh8mDsR+xnDSB+2n9urvbv5Q1Z8hd/IVtROfRRJfMQNVA7UAMJZvUcz4pKzFlcFnkMEIfAfabb7
ZFF0CiMvvtA7gxY9EIP8Va+kRCIgjcFR+4JhU5w7x9xIGwj47QKnM0d9EeZLP09BgUEI/KKmRys9
VWm3YQfYA2U9GPFSWgPTlW4/aHbMsGWEOrBAtPqgQ58xXwv9rtyKrCcD3NpfUqkpx4+EPjjxjE8t
YddufbhtrmTJUNILmkrO6aYVwYSq2E/C6dO+xBWWwtomdFpy4GHCyaX4/kcOmCEcohEXIuYua2T5
7iehYuHvRH8mNqunKxzqOcC9EQalpjXPZKjCO/lvwHb+pRD3KH+xdeL/M+ovnfxz4+sedo+Zu0h6
n+KvgTZzgNHA6XqWR91rJiCyA41OoW9EXQsgZUOmGzxpEYdRuOTeWP+gkiM/oD54AL1LKUAN570N
MYvyBNTXl3HudJFG817E5tA9BJO+0Fsecyno/FguX6xLPRG7FnY6z5XRzAGLKRGMsUo2wU4dxkg6
lLCIdEOL8DxIBGHrRfLYij9jPW54CuN6seTi20/X6byUNjST97iSn7AVwJcivIPBeOAmLlaf0O/K
gP+5B4QPnHYl3DL2rMHvvzemfnI5+edQ/HqgcwtQQ/YKFhX9rPylTGiTRoprUeDWWM5+8g1p/7G3
MvAQI7H/iqLMp92E2hACxx9z0NG0SHbVPlO4yDJXE3Yg9vVYU6LiMGsWXoUg0uiW8Gl9jO13y90L
nxwLlshxoRkMwYjdEgT6gjq5x4pZouppZhPXEAchcaCsykufszsyWDYWBAsjFb/y13ZmP4zoZERB
TGToKehs2ETt2hYazQMXOgv4xPHkROrtjNS86azZF32ATmJH2ULguuaBzNegXDdK3zBBF+FY+S+o
7bV5FEgR9BTcTtDMOQ/UmIrRBXWVM129C8WU9XNoHlXaw+UUIm13TqK4nDkrR3qWSl84cQjlKiGC
HjsbO5btWPbqr8tesWEkhKDIOkx2Aszp83NOC2gezsFj7RRx2PEgilNrUvAqpi5M+fd+OU3lQM2q
16baFE1AO9QyxCAItTsc49NtRe5WZwTNV42dDPgkBVHwTLlk5ClBXjncGvDp2YYFyayC8yhtA8lw
HHct2uWqLcFO3yPKZsy+8BKHjXf2JBeKDeS4IihI7TA8372YcYJZK5IoXvnVfrfuCr+kDMm13KWm
rmUs4KupXoMEQibyQB6kkrLE+LwL7tnaghTMBSPu/lcG3D6Jn9/a6Rs+/XcOu8Rgi4YMM6XR8rMn
Wt4+8GA3lto3biP16/o6GFj8bFAKO+i4KlDB7vFDnfO3bWhcmj8/KzpUYynsZqB0SI8KieUqOUAp
7DZH/1wVZ4xkG9VwRpJ2E3NALkHG0+DyAVLr6qwkzd/xaNyoy+LuPmiTdMe/9fCTDOYBWOzC3O2F
tSNk0ZkxMLPay4+avNEAKcNv4LfteCLnpoGAiNuHdB9Y8wv9wu2ZoHq5H+pvgrW2xnm4d3PHR/Bd
KJ1GuMMC5XfNZLnl3fYy0FsYaL762MWJMYLH7fFsh2S/BCFev87uEYQhJgvdUrT0rfaiDFQpRqoK
O0Pk14N7hU/EeuzUJzo7uArLPaaxvAiP5Enh0pXV8eLZgj4IVWqyDixXaGXefmV/KWWn2rlZF8sK
cUyD8yYF3AzT0m3QhKnHiX1bbQmgKXbBseaYn2mcvlCTtluxseNaC2KhAch+7juKkUZZiXDmA+z5
gDNSpCmDeOKfnuy50C8EN5cYLg9kXzW0x1U8tpyuqbb7BPgTAeeA9r6ue0pK+N+kTTHyoEaqjnE/
DIueqjdnPeOGPZKrXa//3B8fRg60iriuvH6UvbI+j7neWYtk428G6wW44lknTghN5XKshK45qNM7
jQQHjrCU2Gnuw1PMDRAGIZLl+ftePy12PsL/V6ZvbOz63LJ9pFb3MHDjEStwQO6EtPcRJZkRmf61
RZBGH9pEjhnKAGNR9Bblw+WlvQ1E69lvlp069v2c9+uq2MtzsGph+KrDQf0XTk8KhpchUOIS2MZQ
UJ7uO9kKUbNr/77KmZeddIHS6EpJCTgJuFZVoNnMC6D7J8+k65NZkQ0OSXLECb3zPD7wq+ADKJZu
cCBBQIgHZLFVsvKzT9WQcNAxuAzWnnCTp4brGI4MuwRGnRlA1WGIUkGrUJpWU3uB8BkIZ6SlP7qL
R2fPSXOwAMiXdGxjlEOgT9ITNF2182HAS+DizT4GNeyyLNg6bjBoiOPtGeci8xxpFpHu7ePt+pG+
HI5fZDXndsYDPuzlEcdsOkY4SmBnIPLS7HWFpgIVAdGOUHrU1TBzkA12cqfI015JHwUU6Iin2zX8
LuWqEFFfdqg/y+RWMY8hXMgMT6yeaABCmechfo5W5UGlclrLgBoeOs3vh8fqxU1yBdCQKSLMKpuy
mA/guLbn7xZcEtxl4522zamZCCj7YrL5sQiNzNnarRKj+NmzDutaaDMy8bBJB0Bm9m0fl8uBiWPj
w1dosnwZoK94zC/h6CBGVI0tNZyzfCTik+ZMcr7/H4nVLYleJpNfAiL5mHbrkP27WJe2yC7nm5sJ
z81x1IjN7A3iqlCRA7+soZx0jvzM7Fk1Gni5HDX/o8JLI3iqbiaoWCf0hqMjXxKBm67RpCTOOrKZ
1f0XBxUFlxE9wzZkXGfraUUMcY4TaSxRmez0XH7Jix0ggoscilwwJL7JJaQjkfFe+eHQWxgma9Cb
HDEpkvFKCjYuFyXOdEu3VWmzitGO5nKg0z0VCjTJGbaWpCCnAUWHFQt75msC/2lQDCXKxd+GZdML
xsycOYeg+78AVoYNX/LyVVSGQrYNj/qGwBPUDM3Nixe/i8sJTC0IpUrPfGC3M87scuQ+g+9NmeMw
d2yCKMJopTencI4AWYTZKqe4A+b8Knsuf0a7Ri5w+qbyoXafDkMQZWV6MVfylymczBWP5WF46pcM
uf+FvFG6lDETJEqOkAKJNXicPbukqwLzj6Ef3fDS77SA3sFo3WpC522G5NMttKMkZvm1p+FV2tE7
vVhS+0h+0VKUimBZtJEEseT1PSxU0XjoidQ76oiy0lJrDKbe7KT1xGHVPWtZmRaHpLd1jIqM++o6
pgjK7YcTM/zxYk4lHEe7WL5nXWNuOHx7Z7vQrlpsqc6VMwu4rmTJtsgUaPpv/eOHKOMMSYE2c7kL
VbYX0tHkCM348P7S42hk0xd+GdeT18oTjvV5Zs710EhsSXJjVZNGZMm1Xw3D5qAQZWMsx8rIjVW2
gJsQwy75Wp82zkzLsxUx7O5hchmSmZ9vtBeiJz5pQI3AGxBa4T6DpaTO0qG4VKLiwuD3UOZpYxhN
GUujWu7gsZS6r2iffpJczgCoO4777Lnthq+62X+v2h56rLlMQE41S02NiuSxJ8oRokgz/KBuwIPx
ualQRkTVr7HwqjJS+8htspQqJ1NhtND2fTO+EXBAZqKoqk6+k4/xbHeh982uWXTa5yp0gIdNaZY4
UfaiT96Vlp5tOFD/r8H9FLMO2COn1qMIgkmtuM11kgt5S6lbhOe/v9pB6x7T1oGIZtrQBg/rApMy
nGeT7fzcHrDf3iiPRwgDBCo+eUMTNXk7CYxDT1lGFg1hF+vYMaFXFfj5Cmp2zjfCOYdWb/cGARWk
NHpOZwVKPYX7HDCDxkev9yxFfRB/fbR3nhUL77BNn2TmRcBTMZPvrA3zgFWvngVak4CFHDOonS8x
MCNjpQGSLkg81e0K+k8m2RC6uuoSJbLUKHoDbe0YrJuO7QqoJmq80/6IpWAkJq5FssW83NsXVxSM
Zw6qBgC1zY2Gh5bLH2vTkIMekCTrPuyYAEqP9UHB8OfPX8j/h8MHf/uywSobpB6o7QVm0jxqIF9t
shXcYhnwa5ZrvSbEoeY/oN5ylXQLEj3hG+NM5gwKhXLcwE7+KlASwjrQgbz8wouHZacZc1/mzVBR
mAfS8rVW876UtQzK3hEhZ0i4ZcLS+QUb4zlcBsCnQbrapvWj07ObgNcT0HG1+Auuq9WpVFYcWaIe
AywAYHFnIsvEg4mS1fkooU3yfC6IER3vFw19bV8zSPlK114/mfKLbnEDPTBkuXAQJx7jbpqS7LYe
4GgA1LzF8m7bAOsT9TSXKp14TkmfK55xn9W5rev6g4d9Z682Tsf6Bo0N3mByhvufuGVlN5iss7Ev
KGz5nuHevRL5PWqsT4EutMG+iZsORmShi57tNHHHmHlfwjpwuvZSXEHj9p2Okg+P8jv1afIidrvM
WYjtf+cYc2Crxuy7KUjSLwbY5s8LP2qJBDCmiMsNosQczxTYWbdxLUSwU9vH5GFeGTOrdTGqUIv0
Fad5/dQkLehFMHb6bdva1E/Zbal3qUf4GmNr2kLgXyKgD+1s6ldFKH4ORhU1KJFwHH4DTwPNb1LL
kpF/nRRNMt8zn1zZxS5YZXYxX4RKpRKJUcbGCD3ufn8/o/NsZHIfQWulokBm+4SCBELYCJX3Zt3T
X2IUiWY21uPZAwqTgHJDE9vzTRR2SJt65hzPXae4Tsy4FP9uDMw8mDbEXcv+PfzU5d7KIQqv5RvU
2rlJ0BPdUZkE2QJK1Mdwn4GHVx6luMbAPHHvqzFhQvF6UpiJh+AqdyMZd6mvZr25owo6cWGCQQps
8xgQG13foH+K7CuX3UErT0avwf8yJqHVl3KXgLyJk+lJQSUcH5cU6MP48Tzc5ojuefsWweNHDFfZ
uiuCTT4au1KwwrM6L/mQgw+usGRzNAkc61xowRiOlEneqJ+sdrL4lUEnANffYOMzPoKoQg4uhjlz
CTYNb/tXqrl0pwEFDjEPSs3iOycAx8yNu8V4pISDY8AJr/OhAQkdGv/8ts0gMMIAsTgOiTEgO89D
1rk9fihcn3L+H2o7+5oVBprx3GzjzBhUrE4Un3u7w2G55XQX0OA1mInA+1WsrJiFx4K2Ldwruv2A
hXHFJ4wnOZ+ZAMV/dEmES00OTvT5j3RZXl3zYAPTQ5IjkmVUOr5WcrVnRouVpB7ZSyg+2RTInAl9
+2mUw8VyEY0rnJEZonA+d8QV+sJ9S5aIBpx7oh2Xq2qU99EAEkpMkxxVptXjABW4V+SIYhnND2Gg
0Loi/Y71Yez8kDOLzdgi+mzfUcOmyAHbVdqOYiBBzuCxjD8ndJoEsKWRZzZN9jgve+Mz71LN5DLf
Gk8rfKh4lcFBr9JiFxGrkFTyY98V3gYyQVOf03gicLnFayMMo9cC8XpLqjpKcpklgoSMPLA9Z0xn
HfWKuaOeLBqurkXbjplY+0X3imPeCG6pXol1TU96bwZS4DGP7yacNmMsb+uN66sw6vyiIHOqJwVd
OTB8JG4CMPGrfa4l9yL0vhICg3kfhKP6d63L+cb3LZX5UgBla27lZDeq2LwhZ8IkrJA10K98Y+Im
BSSX7jlGcMq9Led0OhssPIx9VDrDqGTFTYTwsdmAYlFk01yhiVBeTbm/EpM3MT6obXgxRDW1XYzn
ze9T3lkupUKslZcY+ReaY77w9wOqKgkKD6W6MqTCohG/6mELeZg3oTsC8RK7fa1mupHfP5EjXHza
Ia14pwko0qcJZxxBQTX5ObvKMlk612+XNdjWaH7FJ30D8xv1Y/8UdodB6FvUf0hp8h0zXiv6RJna
ZWTNVZIY+EXPJ/3cVUOq7PYYtTGggETgHek4S++4ILxucbLjz8dNRUYxhx7qvf6uevsWTkjljV8G
I/AMjqRroT+pmJ6lrR8O9f5zBQiYCpQ7GoF16X/Z0CbfqLz1eDIKXjgParHhCjxIBznstNw5Hlqp
Wwe/zB+/C8tG/UyzK9GE0mRwQoY25nxv7OQ2CelXxNYjaEy7IfXwaamDpfg3qBcktf8N3Sy2Lkks
GU3IG15TmLaw+ofuVHY8lqct9H7AplNwmrGjId1zYCX4bkPc03BvqYkiFChE9JA311BvbprjTMnz
fM4ElolhDlGu0RNj75Ece6eA2x6XFZaUeYb2QvnjV2OSCTYVhVeZbYWwpiUHP+QuEy6SnnI1r5iZ
LZi7JFgNizktBNjYDCU0RMfHjomYeLtpmt/VhG96BAzOrYt6dKe/C3SDAjQEik/shlnC3hwYe8Ai
tKxQ75WuThmZROCKL/M/KBgzJvP6rbQ8ZOVTFslX7urtwVN4MeMmFRbUajH2nQoKagUY+ChS1Qd8
s2krXBDbE1VSutl7iP14huJXRw3cSkntVURw94gSVaid39sZlGQnhzWWvfTIodjZPyTZ4NKifFq1
vyMQMrFkk5Fr1v7+NWt9adLAdXnNefBvhUxTWYb4d5T782gaZw6O12jpi7dRlk+EHvqdbGiW4zJF
NOaxwjeXzJ8cz8pxa0/ApfudnNjkvWtH14I0OU0m4PM7uA2oZQfovHGO2U4X3hqXeO24ufcz33wi
pWNwFp6y1ngvUOY1mHBHJ3EuizsNmdyZqU8sPxf3G+srWqfvrx/5b7JDsASgniWl/4A3G1DXZhpe
2+B8IfRri767AoJdJ0hteIXwIxN10V1bObzRj6wipgtuuVCLjOh90MaYue4QUbgGiY8lWzfDQPUC
VaIXNxfiKuCBWsgEj3HQU20stNTEQ4mtpnmQ4chpRFlhYDi5vQN9Rk/kChWKTmnfbyyQicLElk0W
gNhFnIbvRfV08t6aUd+SQZotMjrNnR9zbYm2b9gmEWkwUGPAsOZ0Pt8udgmwjlpheM8MqspnTPaa
TjrwHwfF+lh9i4qSJdMv6QoE4fpvjWRe2RNwQgEY80qkXkoqJEC130NAnnIx5WV+Mc3gJaVmZu0W
oLUcvpF+bkWzZG4r7EQjQheTKFtY5kghF/YlvnOnaGtPa0ik9vuitEU7If1iLLcvXn/5FpbhOT4Z
WX6rcO0iKmEVZgcVIFIX99XBppD31x5xgag0YyOQj9mEO0g0hP+NUWuyiNedcxGEacAwK4bmaE9Y
i7mF1LOj9leIivcPM05VQ74WnReWboVC9vBWtfFVEWZhhW6KaHxJOIm8sY8OMxWKHla/rBdu31QN
GXfdYVrjKv/Gsxmi0vGMOobwqt8ExaFbwbL7YhhVviiVwMwdmxPh4a9TQgbGfPzUF3jWtTqBDcLf
EsgwFouf1QJlZPCKaaLKr7YX8X+QhxfiZc+OF3RaJEcsANyAtxqYKViff8I4trr9RHYUFPhPpLoc
ZG56B32U1w6HSmwEuhb0Nalek6P4ryD1kM8fA/19xuo3HcCv7Z29gXCEfbeAtNJstm5zSpK9wFSf
DdOuggEM6sHbGosqXCUoyUlNXLa0XHXpbtXahF5OX00sNhgrTOhJKj60HMA7YdzZW91cSordHIwu
ULzv1hw1vkjM5BS9RhrjJOq734rHKRJoZ87EuqV3xPp1FhCyXpZHZ2kXWFnTmAIuRK4POoiBnSEv
Hr6AvyNzcNxUoz/v7kPaRJKmSIJX3bXJR+7OsUqf+aloFkPprmb93QgRZsA4/gk/T6+lxSbhFrw9
umiG/bNhiFTWzhRshU0HwXRvpr/ETp9d2GpPT+xxSYsFNDEMcv1kPd501zjYIrXBLBFAAbps27US
eThn9kb+C6OzNeupWlAV1SMwM0vXMq4OMGEhjugFETfE6RQiZP9NhKQozORCE8XIdO0OJhQTW8gQ
uv6ZFiOraVhXD+EU5CT/G4jBQR2V6oqVsrR54BMV6/O3vGthTG/oy6emFivOLAEvfBguQE8zI/C3
Axk3fOVwft+mUf4leLcvPlJzKm43Ow3FWH/hqLMjiPGQLZTnj2nMXdzIceNrwIIiw3Z8f9vK504O
tXmmMhKVeisn5E6I+kiwo31/E9mE9ttA2EYUkUxot4M6L3uQXAUEwlnJPksRH1HOrqw9NNOKyRAh
EVibNvqjFe/YaYKiktqwpR0VIGGA9QbOGOHKSgaC9z5zY6hfl6EtCoIsHfl5wnmx0xPOCiP+OZCS
GIk3BNVBPYahxOlATXZC3BtjG3w4cT0hv/SnzVr6xFmSxd8blcQuIgAESvF+atghBU+5V5wgc+Sg
1IORezBN2lSrqUiuwZQU9/1IkreJ+JseeraIZFcuuvO+vqvgoE+rcyMiacw2UQ1L1Smd5KpGgGD6
0iJXOhkRUFLdKHuvc0C/5e66BdlvQ00vCNsIFTQi0s6yikBc+WEYqz/HlbZixcT9freeHblmfsFi
MyljCaJ7vfpH8o9blpdOs2meQtvf9V5gWkEKZSXW4HJhLvqvohmJBcI8RGjNlGS/yxKLUK9U7dDQ
bTGX79tjo2n9ZSbWfYgOzgQ73KWr1JqosSX1ri+YoakkOpcbS+X4aQw5YpcBdB+bFNLYQX/MHTZ4
6yS4t738cbsrhp4WJMCNvCT/zjyVcQ7QJ2NBeU88FxA7GfbE/HcE+BNb9hPg9reh5TSCJRuNtZGl
82Hb3ZUgJu0hqmzK+H6xqWU46IGql51ny2seyYxhlvM0VmlkKeqPUoHaNPHSR4eVU1scxHBSTYuD
DIHHVRX9yYoUckq3KuLZa2rqCvRLcE77BTDGaJLQ8TbcvRW0sIHoekH+ACPjRSFMue2Bfg2f2Jra
17WUhgj5vQVD4Hsva8pYoUd1Ura/lKtYdwxSvPcZTXAqKfTGCWkTjB8HioCshZL1M4nUmHpYU+Bk
FjBnPewngdtiVdrmOPJXqL0NIzHtO5EvPvRiJfMwb3X2YaRfjiYH9G5DkK6JF69/jlv3kGG2xmL3
yP7/x7KdpUmGR6QgDhNtB5qcv7RMBBrhcWDvApuV2r40wE+jt+/eVpYAOoBotbZd0Z1EYzKJGXP0
Zov9MbaBx3aKN0Ij1flkOwP8tG3BJ9cfc4TZdnIm7Yb7oCi1kdMgMER8XDL5mcw9znkYXBDeczRn
PUOf5b5pAHFvIYD6ZVRFibnFVP8QZN2bKwH20FOFISNmwmxJb1s9zKB8Bt9t8bGaCGSgISGDbzOM
aF9kGtciDaQk4vQBye5NfQHL6s20eaYWXD7fbo+Ze/HHboOFcqQssGmCtfim4kKs/2s1IM4BEsrA
ix4TrVAOZ2UdYwPdI3x3guEnt5GOayo3r0Ap0LXlAbi1Vpku10zUNfqRLb6x47bqgYm+F2ot3/aJ
jAB8MLnJJrKbkmdxQzh2wawXiDuvSKUs1JsF6DJBSFrmemTWHmoZi+QC6BKPylVDvkY7xfOfSMIZ
H3tT5jpul1W68nSmk2FezVwAPwyh5JHJBeUj4N09jgf6Wpcgon2biEROGIcxsm53djeOR4ivHLAQ
PyzSC/KY0zzSMMndL2y/dOeegutZUKTliSTnTfIA2LcP7vAl8+Uhtspn7GO8QS2WcDgkFNtHWSc+
fIIaJafeUHihGUn839IuvENoL6qwqkKk1cIGHn4uko3sFyxH7at2u5tiCR5NX796iy+xH/gzYow8
s3zLyvXxcnC80KGPFxRE5CEO62XWIUxrJiDwpUSV+rD8bCVkyGnerwMT1h0nn1AAnYf+wnugJSee
wWZ7vOqRMlWrmYVUypgc4A8W2FPKRvQnyEflxALtNO9fTdthD8MhORe88rbmpsHro/7zyBLOqTmb
xRfSG4zf4j8Eic1E06FBNBpISNrVyC+qMEk7OaQSW6ZFDOy5AfZS0QF6PIqpbr37e0NvzeId9PNR
pca3ZtHeXNuMbOwhflGuppApAdU+cHoLwmG/sjLJtoYG9lM4X+1U3R3yYd+RD4PuVjohMGi9aXun
a2/BSBYoBJu4wNf7zpQLZafkYF6FbTqKmIhlQzQOenA5uk91gcwxE7GcHY8TQk5Ht1BgekDhv97m
dHXjSSmLQfaQdEgcDywTqNLwPMNHMpjHkg13v94NJ79uauz4PSVphvgu8t/T6vNknMITYZuVeWxF
8NqWDQGS42HH6nRySVW4oGwwDrBtPzJtChOwirOzPjLkuSC8gX0Xm1/SVAt8LLPxolXdDrHn9n1L
o8Qrug3NTUwTF8Dw5eM8+8ylD7W5+js315fgC/UgusqUJyIma1s1sBGB6gBnnGcEUik/HoZx1eRg
o4naE6KgW203fotolB/U27n3zy4IKe5ZADB/Zn5SyogaAR3fJcKenQ5tSIJ76iVKbsAwxJ1jROQY
WpjrUhZ6VepC8vmTYQSLbO7Vntkr107wTfxSIRXpO05qqmXJZljx6/2fVFCSBy6f3hVTF1O4G00x
lAmVOAlUmADyviomsUfEXsKfeNKAJi5+x4ultB5b0IqaExjQowatcYgcGrv42beZvPjXWMcJVq4Z
Wb5DCMivESzJIW8YygyAP76ZL4S1mthGbtDxFw9H5QDjXSEWy415Uq+XOr9PuVSQTM7OgGgu+wQm
vhZUjJSLj4SLQFZeM7Y13jZz9EzxonitC08NSy5nmCgMiwDzFRkcMR96rmEP1nkRixFvA6GZEIqr
ML5dWjv26WIuux3Gd4fEB67On/chnkvT5W/s+2J0c8rO/yCNEpSHdeM+bdmoOIbWAPQfJ733C6XD
vPfBU7uJwu6Q2JruywZMaedOJPxMj0v38gswSph8ymiR53U+FVSr/1A/rxDivN4w1nl9dp/j7YUp
sLRH6wMLY1LArqGAkHdmAWIWii9VZdjU72eq671W9WzLLV4hAt/N72Pm8DmMxZwqXnZW+KKbVtls
5QnJN8xAoQFwz4iT8Po08pnPEcPnGPDY6YOUWQpXkEAsRIWWVh+hyn4z+bPS8RcRCHy6orl6B1T0
SOn+tOlHo3ENl887esdckaZDRamwj5gtQTraI53mBOqUd5OeXYyTujR20krNRALPZxoXwiijTlZ0
t5KxIEXHJ9K5VSiHWvHkrq2s/pJm6fOS6APuitKW/n7DtBl7OAQvB3DqJaNGI7pBSsYBbphOVI3o
MKaF/b19GF+lgYxzua5yiYS5+xuc0grqauN4qA5joQ1WKboRqE0Deu3V3EfRTLuD3r6WJdLB6srU
jdBtigJkU9V7d5iL3uMNO8XZewy2gzPEtqJ8KzcT23FrYJw4nPc1t2tqhOs8qYh1OMiZaI4NJDxl
WIfH31EZRW/VRuTSBqLlASZ5A0tdjrPMIcuwgET6fT2bLotsCPb93utARai+KRb+p+3aW4ER2GAI
vNTUr3yqKzI7ghWK3EykvNSGBaRdgIZtxI5quRKVb/hEflw7hkKM6kIhxFFUWn+DzihX5GJUAKwp
qezprUjdoVl8Ki1QAi09zBirGY4s7xF0BW7iBcsWlr9cVIiNrbJ7f9ejICjT3Znyxwq5FLA6LNKd
Tvi8Ofp6l85nw4U+DZYC+FWvoUTJmhegWWwo0EnjHo/Oo6CkrKvFhlGZ4RrSXl/IXXqZ4ujMbQlL
d29U6WPkpgAbLnOApEYbtniLWJTAbdck4nNJqe6rNEO5vZatb82pOD68ZP6bCM6bGak+8/k+74mM
qELHrqT+9J/0HSW6S6uv02PF3BIk9VyWJlrkwDzCbq+iKqpZCGia3t/Q7Kl1BO94TPCg0dcsqXPW
GamAnZQ9ecbRlvjtvEuL8P8TtRz9NfmCdooDKfgKrHdyKbsmMGKwTQqGCnMxy+gVEcgtgdqGaXRQ
2M9fGLzuxCwVCTRwozwv5M9nY2Dh3PIsFm4f2eCs6FPpkbziWaf/HJJ9qvR1BzkG0dYn4v26XHuH
zwnR6E63TGvLdnv0dCWFGa9EUzDrgremDA8MUS8CsxUdD5pYdK8puxVWXlT1qFnyA7BkBR4Ndmxk
ZewOmCqQ2FY94Bf+e5JEmPIKiEJ1c1ccpluCZiQvjS9BTmWqQySivjI75XRh1gtRbSi90SNA53fr
giRHJsBahsloJj6LNhI4yVyvdKlt/H8gaNW4xCufsjZ+yOxZ+drriFSxRjeQsP2zmpIYLVKa5gdx
SOubqnpG+IkHtxeykh/liGl/XnD8McZxkXb0sp15AN/+FBJ8ozp8gwjwQ4vuQJlBSFlv0H0GFqbc
LNAf5Ztr7OsSUXzH+P9CR3KDRaKYORNWx3q9fExfgTtLI7YEReid/7Lie3Stfj8MYEivVwq2Hv7K
7x+YALloSEZu/Mro3Z2+kSSkTDmW6ASKQhkwSMF8P8GhS1Xi4CHnUwRyT+WtyYM3HdVgfYpMPVIx
2LAFbgW8PPpC/a+nwHuL2aEbvJl/is5IEiobZGAuv7vMzh20yg/eguOTi7m9i75X+aAveSD5zCek
/eB6XzVABsi/eLQfOs9ywRxX1wYG+cvEM4XM+eV2A3A7MaZ8O/CwG2+hZlXJZNlkRNh9qulzf+zb
28bVrBQtF7fGfrNZ30ksaAmPGC0A0rwrXP3SIuXIyiN/T1f9JnJ8NUJtoX+ZWH3/jmXuMR3q6vXe
oZwg1l9U3IXIGh5fl9N5WaHPrktk6M1jo//mml2etlxbgQSXBh4ySu1Yla1mNYCf7eVLv7gyhjqc
5eKpJaFtHBzKr/3C7Nwqpr5y7Gj+szOdjWL8wa9hDNN0s4jR5WANQb0fju0VT2r+6PqiqLArpe4K
lN2leKOv803pflQljqglNaPAYUIk/RVf44SelQNSMORvs1oUO4BAReXY3nMSBkR0tmV/ynKSwiwS
oJ1DlKQhfHY4MrI4ozfOwgwDEgH8CvwbI5uLe1KVoL4yBd2fEKVDxUf1Cy5x6A157PD0lJ5gKKoW
u5nyF+N8uymI7hRy+RNB84+pjsO+jCLu1Medu2NuNh/UDMOKDk/4dQMmgoiU+6dQp9Fo1pIinZo5
8RWGtyHTEBSFERcqYne6EJLbWUWtRkODaaC+dSPd0YIO2lZB7D3sx7QIfpFqUJz6JabYIFGhdO5t
ZqHyUfio+FQJ56BMEpeYV0jGL5mj90Mrl6eXMV+GlZkLqW3rjJd6mdZ3lx52dinS4XyqJT/guFoo
0MjM4ephrjLbd1g7qNGnj9l3QYD2BuIjxdVc7BqzhdIfmUD8GfAWwwmBrXf4UbKqp2Iem0NkHlvL
YAtu/sQLLesp09WYMaQO+ApLhtb0utpYv9FtnNzClXMj6LPYJChz/I5RKLZzMCsIImtWE5a578SH
CNEZUydAh6wmcCzXAuGJ8kmdOH5DB25aknSzriQB2VTxITEP9F6+I0z59bKQzX19LHT5XJ6LvaCh
80zjSB7BM0onP42AkVIdxIQYtqCeF3QedDUPPuuFmwIznt3499LVITaYy+U3u+ZI6VrmZXDGwENu
g+3+bQ3hC+unBOwYwnjtKtVeV95DQr+L8y2kJhcKrSjy2YDbhd/jCOno6YEc9TjK1w1XTiOqeDwS
e3bogesGtBwCzWyxOqSXL052VsChnv9sNL5evjh9bu8Fo/K2x0hNaLKnHqFC2bCCzCT3JgbFmFkx
oSrX5Ijo1mNJu5Ei/5JVDZriR6cNzYNViiSkQ7s6CD4c3QaU2MHkqxm6FhwFAU8BN+LUhW/ZYOxv
CDqmGPdGbuBuWpvT97ze7+Kqi8FsxyNHvC5BJD3F/7Caht3nf6EhiJFvJ9aZya4i8bYuTALVfvBe
hV+gXCUErbb0xqWS9z9llzb+Bwe+ZTKuhrQKWNNQ7gSg3ZY44FpT64S0faRqURSgaHboUBYscB//
megL2XMmscSKf3pfCSlVzfN8VrneGQhpwwWQxVTQMQc3IeMYjt51rTWWqgaxS+EAhebPjsw0h6RR
/b84qPi02aGI+ym3gCoKcj+mAx4Q6grbnv8k191Hz8A+hvTfMG4wPs0WDdcp524KjG8qjWBCpoMy
Ch2DhT4QhDwYy2T4fBQDrY92VfbFaOg3Rlog9VTuTYbSlVHgjFVg22fs/p8tYRj/OIeulq8OJO0u
q7sDpysBxcx60gQBnJtdqoYjFY23BJG/i5rMVQvBI5rHcmWD0vyvYiVXlUZgvBqOCVo5SnqRgG3k
TDw9eHb20PnoRMAnM29deIdcxJf540vPijljJpOTk0mFh6BjBLrJgmGRSKXznjUEsTV54AGszhyi
v3P7dulYTcVUJ2TTYH4PsMK2EN4H8Xqx684nCZJZi/Vi0gJJ1o1GOgh85Gii/YWAiVT5rpDwyKUI
xZBI20YkHdM+4PK8BcDctoi1MkzNLhBMZk/anOQYnuxrMMzU9i8CWcyN719eurhh1WR0YoF61Z8O
j3w9Hr2GSOX44P9pI9vJRD3Zj3IPhfd5Bu6KexlbncrCxL5tzXiy1kKp6OkPtYjpOrn7dkuwnprf
P9Hkinc1S/BV1yTqIf51oLBXH8AY4qV+tAmc/7EATj0RMp3qHonhBwrCCJFEr9vZSY7j1HfMKWhC
T4gIoPjsEio1VEp9xXfDsuUd6/0D/zECoXSrbo09XIMLAXxdwFFm6dSY6kM0ziY/Pc7bLQ+3j3Q3
/Gim1tHJ8zW1AC0Q5rbN6sVOiEfbGNY3kFAKckW8+YSRNNGE4QNbo58GTaT8uFC2qkK7bWihHJPv
56kDex/4yuNa8IlJPvRUTmUk6hn6c402zChnVp/zyAe4zTew7ocXsJXusO0mN5AP6OtAfe+NzVK3
6KONu6PFYzRhf08LO50h6uLKDlTHPgSwOoAzT+Z7HX00g6jAP1tIKEvKNeBzi3NEiYtcOrmhEEOm
P65ki2+EPMA4CBeKWUuMLTdskZHxZPEOYhQQv1Hce4guGA9ltfcW1uNYsobtbL1UvFmK6kmX2tQd
QuopHwm9NIdkqlb2nybE4fTUmtdKcShVEjlXn6p/LJZJ596uerxX6ivBrQCeG3F7eDmDfac/xK0r
VT1IDsE8pouso34Zna8tQE9fgv8J67yDVYmPay+vH5PVQ/zx7UnXVVcDacPl0KKjB6DC8E7dHsED
DiczWDF1lSjxH6G2BtooKbTadF2erHBoy56SK1hjBTky1L1DFvKaeH/neSnWAcEIMT2jajifETSR
+ZqruimPg9gQzcqQRakUMkLcpUmXn4caOspPfSCNuw5qiSt5lrfkoXF89gIpg0FNmgKzH+ifDU4q
K2bicad5hDQVt+nCB5FXm8Fp7acS5JGm2dyoR2Lkv8hLjZ8e1wRWBkngt6qMOd6Op4/RisZVRtBM
5rmUKsGy5g/uwIPzwyNX8p8qs1OvQM5yrsyyuix5klYQJhqGQG2wQFh9BtvQtjACHoyW4Sz/xJom
Ibx5GGTB2nkhaYwqc0qBTRz+FONKoO+iIbUYNx/K+y2k0tN2Z5wWVI3IZkD0V2aqoBZiwvq02ewf
XDampgBiIx/EHDoYdUSW+3UNMluJS5EjqWh4uW9Vg6cYnmp2ChO/qcO/l4pki2dfnBMe4JTjJ6r+
Nz2QJQOPMubDcSBnhpl7Bk+iPsCgP+GY9yMBTgQfbp7sTq+cJKcyLiQ8WOUD0+9X+9sqC0LIaVvt
HlwmhfFHBjGMRB9GRGilOaaSyvENnwdYCdaSRK2E2Ya+yKmhDiH+JEhXmBqZJI60MwDuwR7zAGay
qZ+qw9k/WrQkbminUEn8lpKVxLsrEj4am8IruSDD1q533zeSmKkx9iafD1CLWk4VDorrL5FxffTc
fDTxW4Mh5inQnTlYZu+p3PLkuzHqOYJFv9Jq5gfFWWiKtMef6RBLpyGfbctUm4+RNjui1tDOcPqx
ZB6fSqp/pyzaO+YjnRzZVYdhy/A1GiWt47/Jn8/UyC7Vx5G+ig6G2wTOQFpzMkUNnxOx6BQcfupH
w3IBTXf6+B7hyuC8ISv58wCL+iZj3zhrYmsLtKL9pIkPZ6QDB5bb4ywUXfoffpY8/qhm6dEWXVT6
QZ//hEHuVSTIVv1fMZNJgaFet6QTdxgYMcqQuEJ4/PK0BmWkkQdF3W/x8AXZUbeQRDAcuJE8vAkN
r68+msJip5vclVd3wpcUsZPCTuG9lypD8t4d7BwWremwOnu06ilgkdyHdUT2ZOIH7teHzbbdsDf4
8PKpp2KgEAvjeUUXfdGfc7v7bAn+Q8yHqhHHFI+0xXu5wqMsY0jDbJiFVzi9WD+0yGP6jS10R/rk
DVNNeW87vysey0DIciX7niie2TR1mrfJJOdSoLkoXUIF/vn0GG0K7l/SENkT2kMrG6v/rUTwU+F3
jfyehLrJ2gTqLwW5aYmKlyhLY5Byvrjc2yn6k1yfgFb+RHLpPZ1+nsDrw6uQvFF2u/k6/nZZJ+2/
2ox4tcyf2ms52XJB0diBfwcUpc2KGLJSxFI037mfzSEaYAgumswu+zyQTmVBQWSN3GwsbQsGTGLB
NLD9VszuV2JTLBMFuR4ZjfdaUAGCK1Yort+PsDgpGYzOJ+zcQFjGWWR8qZwQdYcZGUh5ajPyTT4/
ao7n97QKih1s/R01nmolcukdaW/YP4Xs48aqQdFFsU+xZSMBlnsxZTBOmZDkqiAwrBW8j9DcHGe0
DIkdIdlNC8H7Fhc7Q1kwF0e+uqOnYMNPoal7RcL/4xrKWOaVwvSAoM3O67JaBFrsxkCxaFi6e5n3
mkhEY74xJs1nk6OoCmbylpIn8q3bosl1DoCkZ47NQhUU5vR0MIJppRdDWmZY+4Pti/AL4ciWHY/0
afHI0islDrP3Go2t6WBM4b6sWwypSNqPVMxM5exU5HLehmbbrottdOXRcFHBXUXd9eLYTqqJBrf2
rmZY6iIHxW238YYh8cw78x6GKV9CeQkVULBV/NCoYETWYXzIG/A5/qu69M5Wj0nMFlOMU1q9AKjg
3Juiav4Y+OKA3TbBSBQW43IrA9tHmeJFGlHBk9xvM4tXN5EweUTlawM8mM4AoyYZDeNNOIsruI0u
vGOPOpMfhqLHemWWsQ6/vue24W98WB+Dq/pnAJxMGHcRhjosFd8FJmmBIQ3l6O/ZVojAuy7oi9zI
ZTW/YpkjvRNK6qiIHRosYJlCnK/zpUk97cdXNNIfmhVAw4nJmTbTir5SwBSCb2Up5P0vjOVW6OEv
CCBTfuM5XAzj3S3W8jLwEcOrw/lhLDvO7FuIYBrwYt5eQFHH7/WUyfBvJZ3OtliF9Pms9TsbPH9h
TmsPDWWO87ne0zMryFi+C5kfnFO4qWf1S5bskbxHpNzBgoodvYq408/CtikvnKLae7b75S7zw61G
sfjsDvPG7ZktvzC4Gwn3P4Mp5RqEEwPZSlQ7XGa4f0LFZHO/Kb7yDlvXA/caI500zVETS0nORfXe
+FHofgaP1OTzC5IwRc4eGY56i75GBJy4j+6j4ZV1M3/Eypy/Jij0p9aqQbCKt/9/xLOUoCL21QdY
3kcZeEDL6Yb2tNXNWT5pHOqt2Buczfl1To0GgXUI/Egj5n+9PaQN9AK91xtN8kWaAJm359qBfkY9
wKLBG63Z8dukUAStpwclZHxgtWYJpykt/+VOw1jPWTsdXtTWzLyEFdpCm/6W2AJwnh2YoznCufUu
U7JJ5k9TjAws0dL8IG2ndYqMFTIFhYLWeBTkwdzVnMfYe6rcOqmAAQqScJQOnCiX8Kk/7GilT0h2
/yDgQixypQOjUr0b551v1EcedGKgy7m/kc06+6m+hqyacWvhq3T8N/ZiQ2h9V51AyMUZI4MtBa0I
mZM9j2kdSWlNhSCazx6+2r3iVB5qhKYdcnKH1KfayBBFGDjOEVTxx6h0UEC5yCvOCQHWUswTS3zy
dPQNJFQSM5qSKXTJ7xickPyGXnbO/8EYEY3hMC031ka9UojwQJWgu4xBHZhaabnTJRlcq8mO3YDk
V/q9G3QxS138Rl2wrQ+ryBScIiyBfYxbOHx4Bvl9H5rCEnxxLb/CVp+BxBuJf45m4hSqmd4t3EK+
rdFQGkxRzUFQmG44SGDTd1U0m0k3sizie7BwzlOInMh7ZRfcHUL0nwc2FjvnxQFVaBJ7dkznHkGp
T6hXfz/9qWL8cxB7smLz0AWS1VEa2VbC5Mn6uUbEqjtO60bsezZN0YEjYJe1Ate18ySnLrkRLYKU
LaybvMXgVnMEQYhTx2tm0LZasDev3qaRCOtKCTZcpU92+PkfzbJg3/GcFM1CcbZh/LPaenQ+7L3J
ew1Fhc14InfSzwawHgj5LKOVtV/+5M3QgVHIVuAA8TpinovhHraIdzrIcD941AgHsX9gpdcQpiR7
s/+H+H6X7jU3XUxPdxczdFh2KuoF5XB9r/361ldq4qZKqJ6O35zbOSu5pc1R89F1kBbqI+ZyRgKJ
pr5ydB8DZbFyubqWKYr+XxjEvkmG5+lnk1UxKi2cgaX3SmHVk0yYliGHNrFTzW878BqbGALaf/bk
NONYdde4VPZtgvkVY6wOa6Q73x1VgY4mDe7Vf20ZmdSwjdqOWdhlw6hKECeIBvedcTSARe+/MhKO
iC75hpGMmYAn9ahENLOgk+VLwu+UM84Yyjme5hSVDwtF3tIVu6NOIZZHRHid7auWdFikm6iVanxv
NZA020QtRE3hqcfLV76urqckF2Kue+mZZbyITKExCTqAhEOZRnTQ4r0apNdg5EKe+i0bKSPmQGcW
RFg6uzhQfctdCY7LN2mOu4yDJCc4rP8Zyd8HPRqDZjIYPJ/8zE5wHA/HzYz7OyjA3XTG/a/ck053
crzBL32nlCnnfZc+uluhQqAW46GBm0yZslLXoIl2Q8z9CxRMxt7yEOxuumLf5PrkhDYhtWXeahE9
E6LuihKbLFRaeVND5H6N5F++f9+iPmAIjWmt3OtrRyZlDqDMwP1jaamEcOalzVUr55UNVBS3BdDt
h0XWvzpB7y0bHs1MPkMexBlVvNZhrICWc94Fa0V4z2aEUaBSAfFtjVua0Ak0hgPbTTgRFq72vFSr
zwLjUTXEFqSK3d43I5f1i5+rm/GNNk6WveXjYh0JftgRgEQhzdxfPaJFCKHGHFohEQVSXUh++MZT
8sLkJKkmHD7a9BTGf16mAEPpcYldcpZDI3ubEH2J2glc+ZWB+v12HVpY5EqkGoKT4wnzBOY6m1K9
KdQNnBmLGLPF90u15Tnr/dCrMLc1coc+PxYY+fZ167mfBe21rdfu/Epm2CT/5g0BrsYjZrP8ET1/
tdNIBx9VJzZiW9TwS3ilVFOJRKc3XlUI5CYAuy/H38qVQuW1Vc1O44ZFMDODnuN9MV4XMD5IBgaP
7x3fAM+5ejy3nSoW581ARFRyycxfkCK9NYpcgyFTtYKLgyEO+EqinR9QeufFf6n7m0h35pF/LkT0
q8VSDKdrj7stnZSUbW812EFB3lUTXLv2/+AHCBpLi7dniI6v6Nncdx5cDVDQGLMLmgkT5KFHfj6j
4YTsbFKeFp4k13u0PrFBe8Y8D80oX0k40mnypUG78son0TB8KELWWokV1cW68vm0aPmsMRKdjI6I
GIuO7Dlw0LkGeI+aoH84AwGaxoSfeRYWCdq8oa8Uob6Y+ubMy686jw4AgbknR55+Hkvpx9Q8WcQa
XH+WDmlAP0WJTurjktzl49iTu1Qyz0+gCiqLWdLyrR5Hzf0rMHDXjkZVM6NzalIqFNnI+0uJnA2f
n46yTN8DY6O4Y22CfhYatN1FAnXJZeIFJdmW6EQMJL/tacUQTFehEVWGOnoKcBlXaglX6SWVcBX1
f5eC4FqkMTtXHBGQkJpzAOSDFClankUrB4FHTReBVte9NYYO6MSSKXxDoCc97IxktszSKDVLDbin
rL7691HdVKGr6t6IUNzdTn0MRz060Gg4K4LREHGW+UmNThhBjUslpPfi1Z1HM+QHkw/35ToIhcHQ
ThYedgYNysExuPzdppvZlFywpt7vI4gLCzbIA/yKIa2FKITvO8u/BdDZqdId/RL1NI7VsZz6dE52
8mr13CeQYoqjBuBFWwuDKL1Kd7w3FwgmdSvZZ0JsX7M8Ai9x6cG66XNR4W3pDlH54DWvM/sNOJ9t
1RKYo1XtQH2Pc1w8emPPvdb93Mg1V8md5Vv3NduaA+kNEUp5AHNSB23JO1q675CxGfiiRFT/QWcn
zkBgvOwv8Vul/WLu5PhKZOm6iBADH1COb6scXuMKGtnxymiI93YcJz74AW9wKtHAJCTtJwRDW6Dn
6XaJ5cFmFlf493RfKGIJVY1dN8Lp810DmCa0FgerXhKO0Htu0pxpLA+pPyQAxjgI9AtY0ZZbC585
j3JzhPfUvLH72mMVOb5ivLH3ZtoL0N/b9jALzMtnZFNr44HVCF03hxZy9Q9Ch8oKHAF5cudQ6Huw
cIi2fEwU/lkvLtfOw/6pJpN1S9otRs/mzSvEUuLbuEFMBmWwqIQ2VmUsl/x9+cUxfD1JfWx2By+o
jOsSdZoDa6er4gSiXYZZao2shY182RMhoY1chM7JRaczl7Tt/7IYkujBnPuwv6o+ks6yRNZO9xld
2/DefM8be6GlkQ/ETWxyVwdPlen+dTFnzEgi0yN0dpdlgyMAmIls8398MEtJZUzITZZBT/6urv+3
a20sjixGW/4Nc0/Jf4kFg0Lu2yfpoPzZIussGFFg6PbMwrOou7iQojNlRMiCfImNr97HvuJ8ZPXE
8sXsGTtqc0ja9ZVhwDXxin3GBVN5oyqeUNeD0Ei3cla8CLIiQEpxUs13OmDdRYMwseprWovMRwfQ
gMsQpx5OVOr4T1qW8Sqv6Edip6DOu6G37hnKFyzhzS+WYjFxFjs1rjdYjQLRlYroHMC2PclWa1dn
PBZHNXiYRkNVaMgVq+BLX2HphgfXDMfhLiBb5BNBHrBXySiUiRfeYwYCoe421G9J5+XICl6E6JFN
GmjHurYXFIquPMoS+4gpY2jmzWhzpUwzW7LqM6WfbV8QAO/FAWK3oLZiTIovsBC0mdcTZwtAv21u
kFJvDF5buTKem9zNgHO2g0V5LcAfwU/vyF3oi85t+9ghAUiva/RTcOoiXYIMmJFtVS/8B6LY3crk
5pTm0KKZDcOxB1jpQ4itZehUa7MXPPdIW8dR7dfnb1X1FuinEsM1lQ3jhlmiob6XwRTadXTpEzbX
xoEp8WLcWFQYaqyxfbHslsziknaNX4uIYFV4ewf3JnjcgNd4PEbesEdMPxAM1Xf5tEFGRA0u+mrG
enQ+tkLMFvcRydZXZ478INlLaTzqflp4cCteeGayeYcR037BKCiX/J/SUJ2hyzRsQhQR5B3m/xBe
8FxSF7eVyK/7FbGollsTnZeuWyF7EUNbnj7LhoX4r65w8mTdIW5+5v7hR5+8nOis0hoqZ6z9tRCc
ekcaMvN51MrUb8e6DO7bP6hH60LkB5cF9g50cZOjPkauf6quTqs88fszTvO8LMaFWT0hSUsqYvf+
XkSmzVMQRxy82kt2tAkQTCKPLWC1atIs2CThoumtrM9M2sH9mnyaiVPkF4lOdtGDOTXdOGy6BzW+
5XtukZjno0B2Q//ZIvJ28JAfTkhjcn7JWvSa7jJtPfffeCnBNUaAaqFNEB4RAY0aO4xRiWcn7Gw/
3zxZdr8qC9yGDWUgy50w1U5WI18iKpybXY/QAPolV13JU1HJDwXZE/phVNDpGtYvWbidurYO5eUd
jr4izjO09cg1ezRn6PzIL5WGah8mFk4iT4PdFLdI8l/VbbhUDu+jhHcsHDYALy/Td3DQ4S6KLqpG
veq2aBlBk7JQdH4gpiIxpVJT/RlY/wBpTUdGBWzr2CUi2oWrWeQD0JjdkKTb0XOPdK2LlTf9zaDm
ntr323uQGy4uK64Bk5fQLKk4e1fjSPIixbHBIOzKDSZogZomuxLk+QsC7SJOak0tiD2YZTlxi1fF
2vMR1fbdhNX4ajb64JNk79bbBvdcz21VrhkJFx4lHZvOojFMlO1Fl1xWHuKUVhRrEsKU3SpMkMuN
0Vh+Z8z8n9Jfc64ZzgFBhxY5v4meECTysucHi8Tz0c8M//XwkQo6xRub6GFW3OE9mdAK2V22RQKI
uxcYTnlvKQ7TwpPMXBPRVGJ4HjJHKIzR4kRvXcvVhdZ58SETYaMO8tuU6z4AXuBOz8rpiVM9hTyZ
q9dbeZ9fs62WpTqlDDitaqAa4Q+6C5sl0TuFnxB6qaewuX/7DBvA8igS6BdGoU7Du3RMOwSnJ9QW
GsFZ9UP4HplarvRk4Ayuhcaqq4TnZV2Fxatw4eOK5kvifMwNxo1GOsI4rSjsASf7BfUHAEOQA/iD
Ry5ArIbgDJK2YbKrIwJWl+IX76WPy/MLtMn1jrw2nWnF2dB1JbD3a6xzPgzsAd+L7A9A+xSaIuRQ
NmkQgct8hHBabpNLDM1ookh9rPThSjRlJk3EpI9JADwDR4mq+t8o9BmMHQ6empX+/cTYixoiqSDQ
DXqfWTKgJQwC1CnlRdLZxqiypMB59CfUJ5CIurkPviRrzVap8OaHdL09DBXwzMEk3R9GcoK/0fkI
I193KxcfoxUjgfgtLv8TLGAm/Ul8hcVabs4pnw478dqisVvIGBDZewleHBJAKKdr3LabCk7aLiuO
X4JT/Yjzp8dNEbjEz6CBCyUZZK0ZmcR9WazqgKDq9jElj4yz6A42Qs8/KTGuISdo55FU0GqirEQu
fdIdk3TI13rWC8IY1s60HQVRAgUdWXU13aEDLK/5jnfVC3GqHxLKCUugRpyFlLRM1uccqe2XD9sA
tY+PQ4OEF/pDNa4AoEeRUfpNT7XndZZWDdu1IQclllO4aPIVvBFFDbshHj74IkP3ohjA6i5Zb81q
C7yxZqa79hgr0T4mUeCaG6VyRkQpLK1ef5PuRfb5jT/k+qEp/A2xfx8fV9w+QVhKfF+K/IDMyukg
rGrYSoQ0PpM2/Gx0S+22JvYFkZEf8Uovsda1v7skhSNa6GMeHIZI2QjGNVu1NZWE9sPAgZYJRoym
Zw6+U9YeLoQipvIYQBYVQwOYNNv9oY4c/DSTa9gUC6MS0E2/V5rxaIHCgF1YnFvVF3ByGd/HTxKx
r3iWQuzJSDnYesebua3GymAh674yL86pzVO/zUMSDRcrY+YQgeJbqPR+0bLQIeFnXrQuaCLe5ieJ
tYRq53uvqeDABmqjOFvo7bMvydGBxl5ag43jHYhKmn+e37v7XpZVG43jWgKrRArkRRYM7oVcj3Yl
57gEJUgt/7mYaa/jARdleguKVhuMBsfc3OaNC4CE0TehCt7eCpbuhpkYY+wVGKOg7IpmamTkSIcJ
s8o0vqP3R2ME9kCa3lBGtHZinE5icWZ1b6jxkizSKtrxs1EeYie0IgEgbvi7FgwmFYn6BVAfmm8J
6tqyE7/35fO6nL/3aKoxKBqbA8fnCZ+2/ryDlK9LEtLGqNb1MbzCCk8YDDayzGxvKXLrri6pVhhQ
eDfFZ+iOLkLZGKXUldfJfrBK6nVl1cxbtsVe5rd3T7Zg1BusX5l4AtQNZn7JcTDLOdrsJlSCZKoD
kVMs5U3dPIeeif9Fs2SFCiu9Nr1DQdwEEq8nKU2ti3KvxByaPGIa8vQxkN0aDaLaEgwsYB5MVOc2
g9oxz6mD5yTQtwL1n9oZewKahw6UZbzL43q+RihLCQBNiaC6gYf8lW8S62xCbsk2cxEZ7L5Ba/xV
/K4E6b9sEMZdAjihfQ5qxIAgzom+0oR4t90Gew9m6NRRVt9wDeOCwpizoU743v0mzlPBlcys2pRc
lO/fnXNJbYTkFrlW90z//lIHWRdsWT0pB7SznXwfj2mh9pfaLCMHp3AhycN7jBSufdTRXaibQ1ET
3IHHLYxY8UQPs19Xr9sPf+IglGEHYTAL5X6h++GSYUwa622O+SVUqSTej9t9tfmxcW7uIXjVxCyi
jc3engjpKoEtlYY7djsqRlXZpBQMgbgDPERGFIB0h81EXIwOBNHRqtbHX7L9zX0S/bDVSGT2q7dM
hmnG4BDsEWZe1gH4M2hsD7S1SJsMAqGH2eLwwkFKv3oT5ueshTd/x6wpLL6NGnTPVSbHVUQVpfYi
DLGv0Re7K8hjNZDsNz5yvci3eSkcOCX1U1AUvNiyNv/F1czUQYRUqheBFv9TwdXYu8SwjzZhzwqS
ot3VfOAC6rSSS8EwG1/cCOY9f8ycHEkWC+xrTqmmyKIWirnNhm9BmfMNatJM22bZ1TNNd+t0gzAh
t/At1+oQgfTnDzLmNtK7rq5QQa56tX6axcu1iiHmGdToyjVCmiWyMkM3tZ3tTch0vClwDkRP3HiF
4682SrI1fk0p8/Sqg09do+f06vsoEOcljkh4kETVYTp8ddbuEn/Nh59DNJnidQgMHNNy7jXt0paP
iLQbZDnjGFUh3+jiGJtbO6O/DzGaE6PJZHEFeAzBFmWm+7nguNgUZRhFr1/dBhcMNft8MRNX/djf
v/ynJu2Fa8S4XCpsysk6t06Hu8D6jD7pwLuk3Wb9O3bhN5Fc2Btf5F0YZpN+2vfww+OV2KuA0Ah+
hhesS7BzGX19iB9NxkWOSpxNPa1Uu2iGRxWPXgA1IOyeKd3Uv8E4RuV19GOnBrSEmicsQZoqATnz
6fWq8OOGn78Wwvy2EfhHVb+W2/Ov5DoiVeZMsipQl4PUHYItmVchzn31Mz2tO63FW3vobG+5dpFG
MKOUH1NvUV6K694yZsHD0cY0K7a5qW6qAlZGZNp0ma3IrHPVYteLNAYjQywr4N8wYn61d8y6fTwd
OgRRrtKYvT8oJrtMzRxPQ3WKtkx+5h9GzeYqDJO4Ifg9sYH2WMGr9/TeBl6yf7KH57GNW7SNTdRI
TTzTYTrp/qROnjiVLZ4Lt8Uw/yj+wqKT42x6DjX7IWKd19N8uOcmDMbof/5y5BD9IajLT369Ixic
bZ2zFOx3Zt4EDmlxLkH/ssGh9+wqGqWQvcyBtRRhMLhn+j3kjr5Tl2K0JtctKQOg1GeMqPyl25fJ
WcLNtteJ5cX2qV+XaeYPRZ9LwYYJdw+c4Rl0Qc7wQcTAzTcYI1pks7PHqSjOXja7ZhUVST5t7kaO
+UVgvRy70SlEro+r0TBXnNQKjyb2y5Q9Ij4ODFDK3nnrC9QjSzJR3UqLQ19x+9/+N1sb6qtMJXwQ
sjR5cvUYSoSen/VidiTDTyizFK4VPRezQuyc5GZPInxvbytFL7xkRcVDqKRqaL3x7EGXrR+vIh+S
RWNYCRW5Vd4PYv5AgrItP0iVx5E18847bzlQVr7tL+TgH6Wn9D1uPUTZj1mtw0WLPyUuNwGk8Yyb
Kcs9739+M6083eOcEAyO8yfkd2Jg/PU6q2uLrmx4m5P+6jRcnRDRbbns4b+oCaPitKmpBxHnS+7V
0p4iNkZRIeqlIblXjBzK362NoQqKDtBoL93vrBcvGHwm736F1LLYKYF+zwMU5aoMUaURNFwBMN+s
tfT+B7I+f70uBKejXhrWLVlUy1H0uiQW2n4zCfWVi0JPJzYvUgNWqQZ5AkDU/MhsBk2crQAsa8MW
0Za6Y+F34xaMSAit6PXbcxzq28/FkZyQOZ/uPTbmktenIlx3oNJi4WBb+8cNY1nbd8kQlrwzQO9k
eH8O1VQoSDfUEDJvr319OYEtXWQczR7y02IHSEi0mZP2cGpFfdWt/HJbOM5qasn1lrI2LloIHROt
zsUADPfg/jVO3/qQd896ai/DaM1yWKSDHzSQXKc3nbJG8zqTyR6RynSFcv3mp/V86s6IybPv02P5
zcZjXl/i7Vo2iSsfLFLYQxTmW8yFgWUVco8ImdQQ3Gub4DOqaK4PvYOsphxKIfx3F/1U/r10GdQ4
yPP1WpjaCjNBH3UOJ4NCKPfD5mRm4DUg5+9CJ7nmRt+K4fsgxY+ZZs3GidLHdqJp0F2JTgUSI6P+
sAWqVc/UCvGrwQTwbJVLVwXNOQ+82Bx2eFyyGUwn5y7aMZw7217gNa2hD8+SkL7ZybzH1k7xADcw
IiOpddomCOWnJebc06KF4g2UGc5riktuuLavFk5d5GcIkWjSuJ7qxGjrZxfG9/sCJDUFsLWI6p8x
OeB5Iw8Wmd+DLtauaGG2+5mcbhDgMmEP7iIkS5TmxiPA65er8PFuf7e1YhUGoah4a6eaKM7iykr3
qjZHslfPlpYAyC7Hm3QGFTob9e9qQ6Yyo7XyHtlpU2vlKaR8YNeD2KVExOtjuKiKxWGH+V8KZyL/
lN9i8lvkN7NwN/eV3KwMyhIe0vuhfLk6KJ+bxYoPsF9HG3UugZ8YXlQdCgeQDbUcNOg4PDJjUWAb
uTTl52YvuCjgENjagTr8lC2QutLgLKWg9sJy4mzouNGAxzS5j0Hh3wl6AvErVrwsRvb6PYc/M3PR
cXW5KjrTDkj2CGfacKA/9xQfqbQ8eIAsr8//qJDmKAzQ96oyqgdz00gbnRPCrCcZVl5P8qQIwM8f
LudRwZmulcfXacM3IW7W4fnGe2tEBIeAK4tQhC9oxdg7rY9KYbJbUk0sELmh4hgrPcL05cuH9HG9
MoIEtlESf4u5G1cwyaSJn0JZphk17wF5Qyo2KFxmEoJjNB/BtCRZbjuUAP+se0jHNFDoVmdFeRpf
BtXD7uVL3V81chZJYr1NtRYGDzfDmniU5tE2pdPgF3N2tuval1F/kTk/d44nmSXx8KhENlFIvWId
/PBcNAYVEKOjvBS1DznMWN2TSBbENGK2CcjlF+6E5kv5iseUVX6qm8HpZxZVuvHpTxPk9soQoArU
N0y6UcRSLw5ZEAdRcBHjHfFKuySaF19afkNV0UBlfogMiAMrSDAYx5EDFDNOfGBOHY3yoFSM1hxf
PrJXw0ZyeCZ5zGBVWhlj82RQ2DAcs/OVcEq8e7sRCWV2Q6IF+z1l5HMcGptZi/2j/y+154XkXUXD
Q6zIFk5FdpEomP2feH+g+OheDfb+bVLCcRdAbkr+W5dlmr5E/8wy7J95swyCvrYCZRo+zgw/gMZG
R1LI+W0q0W1mTVDmIAAekkv4zm0MZDZuZiCl4Y0e85RHmGzibA+qDtJecX3r8eVbPhLJ0fokRuuM
mV8te5ND/HHjmeb+uRAazadiyjJQuCGnFfBDOD6Lbe24EK6TlfS8DAWvMh5yRcbJ70jNYOc11GwL
YOoGLKtoTf6p0RDN6oEjBZ0rITHtyNwXCHv8JazZMyr0UztKniEbWMc+Onqh+/xbcWg+HXcVWYra
Eab64BB1IvZaquh0g2LqdBxCQYanH5eYqeww6JfuXg7HowgTm4ooHdcjwEt7nom55tGknxlLA0ei
4mMSuhwVbjjEg3zG8g/ZKOM9w63IutNU3C6dKLvFAVJvXm/APmSYZvLtQ0me0/QHXDO5dFXopu63
tYHCzETelWDq0O1cbRyI2OZZIi/ukxFzOuZZCJonydrLA4w4pYRrPOQfn12waLunUiBSb91u3s9i
exNFx4fLC5SO1TVa+O6YxKS8oiSU2EmpoWTW8Po3B7W+iCH0WqFjDaKlLLngu0Vifum1VwtSwno/
/M71f95AIJemNAj0hNacCfuZMBiSV0BlYKAO2aMXjKjv7VCOCZMmfmicimU6skeU+h1ni6k+NBe3
3nVdvFJ6qTMQvzp2EBxbqNYeARVFgZ6qCvrgkWWXkjWUnebV6y3rrZDbpceViUT3KadmYdPkw+kj
Jor+KSJ+jqZN+pK5P/q6m9l9ULMeHRQWcacsZZFdHkruoJJRaWNZwhNOeHKLLgi8HTscw18tA9ue
u1mlE3/y0FA3UvwuR9O7w+7sB2gUMUahxRo2UuJqMlFuoODmGkR1uplF0Zd77tjE+bY/ZWStf8kt
JPzXLFw0ubj/BIao94rcFKzyPBoiLoC6qW+zjmXc6CtqTbOVig4evV8AntGCuXCkkUf5Maeo5FgT
LNtWrXA1qRtBsYJ9z37wLj896wUoaCJaYoTWWR9apr36l06frulL38K5A34z4Did0hSermY9SVCX
MG4nrSyLVR/+PH+BFCchFL6AlSHMBNAjKYaFa8/AZg2Af7G/jWm7ZNDVBxEIUs2GlJTOSqL+rsRh
plGwZ8R3i7JmZo+uWAbVbmckt14nPalXjn0rfbGFOqBQ9WcI/BKeb6xNBkLZbpAxp/E49vN3/Wsq
J8ALm97+UcvKMfIQ5HTnB2stVL9VCV+tAmH1sPViCZ7WfBz2+vog0QaAdVXK2vhYyLqzeMrxiQOO
9w9Bgfiyc+TQkayZOAASO5DC0cayKTFNex2+p7NtGEXqzHeAi4I8alvqdccp0ZiCMZrBj0Dyf1oR
zSVAAitFYYtzFxBUyOhAWBaPodmgdiBczaBtuhpmZQn44Y1cST18uX0LFk9mC63grPVnWgccpUoO
XoTmF+sPFI3YUL2IYeECSaG/+nNM21EsDqxdyAsXNaYm37YV3wIEvR3+/rsL2V6MV3zhGdeZO5nV
whJAYvR9OAqHkp2ut1hNEjW6+N9I1o8cnMr9n7CtzqqA7XIyAlUzCwUfYPHaOnIfbMC1RlUz1MQr
KZQ6EjYMQoDAQ9rLxAFGoktQBuDomMMH9UIVcgE1ZtdUuSbFa/BHOthpNRSwzvZotPMPw4xTL32S
GDtJ8MXewTgwjlZoE5SuGRQeBMXOqTmpLv/wspq01hndK3k3F73gjIiLDAsPB4MM2qTGOfPI8s6J
wdjnWVwcb7r6HyZNJ7CQ82mZFvmdiYexz8xklwJ4VjVHH0rWM9C7AWlSg1T+VAQpK57DdMVOilPY
Dt/uCK2fR6/6Qr+p7sha48DLM13IOF4WMRUscOMJL5iuc9AqtuJHmm1pFM2kyx4qpUVQHT/uPAV+
+3Qf8xxwps6/JtkEhbsDirBcWBO6efyYZZ17HqbmRf2HSw2QrX4f7ET3cwS3iwfwqIr1w/bg1KTU
BUeYzCIR0yVK5MVyt+oAgiJ1NNLser/4dOJERre0xj266k5CmfuHbsPYvCocq7wGuR1/nN2VUwu8
S4SleN6ezDtSh3vIRGhxwZf0IDPtrLD1ZY1GlrTv8xR+rM+vUzSNhS5nk1RKqAotYVUFgNW4CTtI
NNQxG6d51Cu4KP1fd/YwM/1PwXZ+v/LpUMA/EenvtgQBe4mOWBGjnY3Iobd2Pt8EedPqKo5sAsgK
NN3S4wVcO2qWsY6//VjLXZUkHhJJz1cfzwC0loETekELntCKc0KDLn67XLBa1fhCLDKKJEQRKdtf
rN3rD1duA3WZUEn51c1mN+F5vEFYpBqN5BHQYRFw2oL5ju0B4noROhIF0UouShuX7OqGGGOOYtKt
jRKoAR2AAFT0jeEhh3tf3RSWZJfWLdhAlBEBe1ap0x3DV1iH90Vpgtijs2X8d49otYkUaw2fmlTS
aRwBIXlB7pqawWWAwUvCYa1hS2JoRx//MD6NZVtFXmfp6PL+sLs+sO/xZRjki8A51yqKlOKOdDyW
4GH02R4Fn/2inJEtKPHttSCwC5RsIOWDF2l5ANvKu6QReKZIsQSyelmuYTVDikbvaR4TnC7C+wYH
/VU2cWYSef+BOtC16DJOgzcA7UO1FMN2dFpxqkw5A9VLsT/h8b9y03j+/40GGWLWIyuiXCAw8I0t
G98jzDdNJ4Q1KjNLk6ffWUjrbNkQKKXvnZYGrrEMeXtx8MAKw7SgKhfw8MRDVx8+NaZuor8Gvez3
RdEyaH+NrwiklD5oCXaXKDiwTf315KLdBE9hpf9pby4JABnXB+IZaiEZ78INlk4E6uHCNYdHD2HT
FnHMOYuK5YInTuohm/OMwRtiW1JWASTrBJYwGdvdBsHJ0bqRfUexfVDh5CgCacUyFOOzoyHXtWqd
CjEUjkhWFvsTbHVN70fe5J5ltW5Uuj3dhWwohluMV8/rs/wQTonQWkzOKMopk8wrw5BO6y8ccNK5
6oL9RCCjJXq5PVZwz1caOROmml3fNIBDWzXgj//oWjOAAi8oIWN9VcPd4TvX4sujlJDs8HZyGVGE
VP6gCHNEoidtZ/7NNIvmYQq4sCOAixmgci2t+g/iFRsImX6Rb3cxzMxUSCOnlcMSsZ8Hx75/PjuT
bFpOfj7pevdbqL4LnMezBgsmRaiifFDlIiNyLoeb/1y5HRwgIzGqYfufegGj5wwPjoQRwSnsExGg
XGaN9bK4aH8loj2PMVAEuZO4wrNza2ZHMCkt9/optmBHsbWI+f9/lMnHmdzM4JXFczIwxYTJkGxQ
1SGnv48MPvqmBmG0ypzfJuwZ3A9xNhB4Ab02KiI2O+SOOmnt4xfz65UKX0GbZSyhhGOFw64uGexn
gkvrQGQAS/Mdsngs1AQa6KNeaF1WbjafKTjjOgy8BQoLxpcLlJNWnNIEKvQvx2gNO2qOtPUdT83r
djk2YptwJtfp3RW1p6AwwejEzqdENalwN8YQ02drTzeZOsRlMZLk8D+/pNyIGXE6GM7la1n9k3gI
Ya3qLHALrwxvYp+lnHpaQG81Q25+t67XcwsXR1qN52VVNOtyoVbiD3bnXqGtboeSnKdSQTJC2l+O
wI7vJh1MVSXBtp672dyLqnQ3g5i4WZzPgBvsl/WarOOR/qABVFlz+7n9Xjx/bOByN40ZM+i86p5k
zPfxaz6e2T229LZDQszZfMDnHZC3MIg7ECOMhqoLYu1fIaLd32bNI7FFrhQsl+JxjUE8HQdxkYtr
31U5JYO5LNhB1TL9vMA7ohvfGZEFbpURPjCYx+/f3xv5VlhvPXv0jIG1WoxRzNE0mubGKCtZ48UG
hJ4APYJ7A85Bnqf7wgkulzr5ByqBiMEkXJVMFaSNutPVolbBPnoCQUSgUMJFYTA8wmqs1sjioG0z
CMV6kbiIM7shDwZGUub6ZCb8CYvUzvUWE8sDGtuAWgi+z9DP281KqzgfAoMt/aArqDoTSDntb2B2
TEfv6yVne/S80X7JVLqJ42/IHUJ8aeI6C9PPza6Z2NjL/kGJxKEBxO5u5syiocWtp7GsXTtk10TW
DiNy2AEiWPJLTChzxVWf0EG1bAgpnLqUk4s7KC/JeLiIR6JvRnXFrvkcbhKNiihE27eKAKNgDVIi
KmnwDrkqRcKymsV6/yyy1gM3XLVd/CknN8bg02XAkMg/LcfG8R8H17pl9SIYJ8hgb+2xGl2/NG/a
f73bBfl7dimuG9buwooelSn5DlcRPV63t117/ilYmcXUgqUXVy3aawfDEXJKq5CoSYNlsu2z0h3i
PHjqnK/35Qj5zocg9uunsZd8hF3vvLSQDP8AZabkrqAGJJ5ePGALKVZqqhknAdK7v1JWFtKOobRZ
Y/i1TF1BIWCbnDgBvFJIFTUh+WKqaaEXgCNRdgCgGbhx0IKgtJq3LqJbpIMWl7qS2XKLWUmJ/JVI
byANj0nimTS3/7nUqURQCmNmlwQ1GvLzL4aS/H2I3LhRaOnFYAdS9SoP3RPuebZsEDGhJDS1WftV
Eu7wk/3RWLhqUXpzzUXIreJrimFGF0+XBHim36BIodSesPy93IZgKupMh4nR/UtlJIrm7qGQZXE3
w0ROUMVjAsYKj7Ws0UU7zQzUn/uZrv6BlepJT99qecchLSxGEWh7bbA0WNBa3BiudM1ACVC45fWo
Kt8U6WA+LhMNBFeGH0Im7MgQYuABwtens3rYpdT2rl3V9Y52kk2Z4Nwysy8nxVal7CkBUYlzj+XY
Qrp7tDQbELtpjupXj7QzhHJ8zxcD/w+gdKNFxEWiWG95a3YmRNghfsopXLY781hQJ6a9e+lgbQ3y
qfVGCAfJiR3lTHDzMPRELyicLsRm3CdAYtbQLe6azfp3PL30LfF/Z+tgS0HUVlXSK6JZ3fTK4ahg
6Oy2EYoqQbSkQWDRJlqNIRiwTKzzvvG5MAK6mtZakxyqif/hdx8CudTGqhK/gTdZIcWqNQuUAa7F
zDmag77/2fijuhxx9IwQtwc8OG9dqSv8IIuScNQfCxktRFK/ypsGKCiWmVVrR9IpkjcOeuEsVnBZ
DiUxWiZMec5Q6KUHs4oD14x7hVGOrQr7BAJ6qXU6sEM3E2KErlk0+giMcTEaS11CRdiz2z3ijbPc
N/JWVewXHVTS59Ns2iEo29thOfbbc/67VN84U6J7r1QFKcuwYdgPqPcaf47QkbaFusUkrlOpP1B1
xXcPS4RZIILAamcS1HWryK6zb4Nka4ha3u5lCeI4jXx2Ozkre8TYuJzAvB6TcFsbPcLuzXvWTIco
5mmaElDmmQ0/R+kt3nzpH7QYnjdLzpkJJCn1FJPXzgyuHZaiG7D4CmE1dUYR1RUmO1Qf9OkqSRJR
BrzwPTdRCTqdZpXLI/LcwoddFVmXTYzmh0PgeFPBnEvVw151kZT4EU/jCtoHkwJUBByjyIr51NHl
gcPf9Bu/ASrkskY9NkCzAW3JIVPnMAVJDTRWR4/I0bJcoAhBXPBHmHo7OglUFAo9I3dM7q3ui6iB
mS0IEVA+6RONBFPl1ub79PkbxRzowA/vNFqUy9/mipTgR9nDhpB8tLYZwIV4Noj7TLSAI53myUWJ
g2d7hCYt4y9F3RCrUeWc3z+JJ3+dRDj9wXMnSQcNG4zB9CQyxf2TwwM+BUsiK9T/7cD5ssXZG4cM
aC6L6UK9SHTwzmn2WZJS7vuRsdtlwRP98Wl67UtD1VFO3rqS3oR9U09NvMgHsVPEZVxuwhWhRv5A
xX57Ecg6UYt/WLbE4OhbkJ4b3Y0lMetp0AaNe1CucffHUhn45Az9nooU17cBHHLiFVtIRnNJrGuG
Pf5k3WduUoaVnpX4qqnn0qoByfWYWGGMtNH2YRF+if5qxnDe+8g+y7vVJSpdZUdKoEumy7/7AwvD
+n7lpc6PC2Lt3go2zkXNxzuckEi/ulSReta1Qap2wsHvyCjKG4w9KPUdLRix5Hoar0kTMmvuiH+o
xYSAFk3XFjFJTykdbiR7jJLWCqBpj3SWijUwNp2gmWZCpyRGbsrHj4GEOisLszAB3GVuo4QfCP4B
NMw+nQZ8UbJdpRk6QeWISLdKDY8JcoC5C5TDgzfqmO6+WyH/oFxFOikoE3fROmhbylTt1JamxHQw
9AqF0q62aKPbWTRjoeMxIBdxakUfU6vFTdVwWiTDR2q/3w5EA4Sz1lvqsg3z3aCdqXpB+ajMve2a
V/NDsQZDoFnzGm3OdTAeEL2yZQxEzaXSywr5HcRCLIiDWunBfbCchn5lcLZAh/z4LBmeI6D85uyh
6y+9DJXKGnW8LdlpyuIvVhTnAFaODkcYgdmJoknUt6PEBCbntpNzQiM5c5gOItGOjckY75+77lky
scpQi/UJ6BOkrL323l4sw7oyVNkXFkA6yV4u6/kOOl/K+NCyzNuRAjVxHrSzPelwzrV5BMLEUf8k
Q8EDyKh9brOz1RwtPdeIBB5A20pXXoKLvcsuUB76PmYRsqKZhlXYG9sugaKa4rAAsdtAd4icNpEM
iZ5KwsvVYCLdwA+2YVebor+MW5QmJKt567oZ0aPw/buVIGj5yGqpCr5JOakI6Jr3tBLd54ASniJy
fIdretzHBc7cYugvKUJ0CCxyOhK9RcE7s1yqWsYV1Z09cStTBdMm4fpVL5DUmxSwBLZlRPv+gR1t
sZ0+E2nGurZKQgG/ZsKaT6edWGz6auzvsGSsBpgCV5TohoeCVl7LSzZS/0br2k+cUWfqDRM/jH1O
AKU9PCT352q3hF+61YF5RxrlZiEppSLHW20mjfbBEzakxqzbtVKaMkujO39pB+FWKpfqP/7RTgVb
nnOANenCSQXuB0n+/1PfFi9Tahb2LApMhziNW2MMK9XSVUYp367e3Xu1do4JF3mPtzS22G6TEeD+
NPEyVLBdpgOZ0WU24ZR5i2NDPsKyZIoYSUmetN7MNp5ctOpHiBisPFMW+ziIrkRa/R3EKT1er237
ACLUJRnqC0KN8TvrNb2v7bvER99NkDjjIFkHH4e96MZYf9KfVBy5Fu9uam/nLwybkxZxYdlPYPF7
07valbayuBcu1njqCZzFb4Lmc2+Gd1Ui4IrI8RKI0vZrEPv7eT/VlYQ64VqOhx4dVE+EkSVofowS
aetuYTfz/gSrksT3pYkK+qDeCfk/f5ZwMtvuOBFoG5daAMQUKpsChWR84nKfkFv6m2pkZ860+PYW
/dNefNZzYJpR793X4HmeeKXONEXzA9pZJLq+lUHNWGEKLKNeiVpeHeUFHEQMjuS03gdbWnF0P/R1
S8WYSUmeyxYEHs47elN9kJycy4SvLcAVhA+p6cffcPaymkQbz2RVSzEsTSwAtVKfRPkJpZTUHF8F
KpkIJvNbx/ehD+ZhllPaPp2Te4WkD58uB0OdFopHcPZLybchMpvhtXE9JerL1wjthNUc4imgtA3i
vAvLaQ5Wgi0PqJjQbTX6mXTAlhV2CnSIYP/ZeCaobfZN3bzRhi2eoHpOr+hXrVUeAOgq5BaOWVY8
1gncZ3rr0HNknLmnWcV9Vl+vjTFBRYAsJ71RW7/ENrjo/k0MM5ivjamX9p09oUnuADeCYnUaeQ9+
lBW8QmHhvpsVTMyHSyhN+H2cTDOoAp6JV2N5h7SSem9mhAmxVQByIrPKxDiDRENAl68rtwZ2G+Bd
2eGYS2M222yze2UNBxb+OfrTXJ8qGswsreaoRPelwQaouzFU6K36DRJdXWcGx+nfKbtHtFpJcyPT
n8wgR7eiuRyNfVI0veXuHoGImUWfkLW65kD4dIzQVTVGFClrbpEFdLyMn0fGA+rHTzxRiOROQbih
N7+q5i3Y/pWrKhQLAKOnlWRYkNgALznInKRAFYSyGlMd9uWW4R6RFwea1Ny+qDYsTDZCK9GCTACa
4DbTputcvoUmRVDBkVg5tDhS94A5wPPBDPQ1apR21m+zjJKE7t4mD7bQGijAOfDPPhOIxv2Ufa+f
AF5h/7LueH96ICepk4FqDtPoZWkFzhc3D5/Yc6R5ehrxX4qEO96nGLb35t+mI3OiSlCyYegLiEo6
9+fVqfNl5J1LjuxPrwZ0MXwgqDKYwK1CSYdMk7cigESaW9maVUcUIxoxDxSbQDPaaDDzGId9BZsz
3LDU0GAzoysoWy/rLGMzbLYD/VkMzIoExpcXj6ZT2GERRJB1ZCvIqtSeL4krH2SijRgO59cVq6VQ
ZQxtoiiRmgDE/MW4XJa2qKbu+LZO4P+PXFnOrylpPSHXWG8bpD+BvavlA0B4spqj2MFsO4ldUCPL
7UIhj/K8/Nfqo/awNMXI78scA2Beehuw+Rdf9nCxLinbWemuCbQHeFssVtqNb5NkR3LTKQBD11Pd
j08NkRIe3hV7nvu6nZ526XDDjtKZtM2MFdAm+wg53mw29ObYo3oMX6aFCkLvbd21U3LpL5Rqyvd1
DLlETqCFr104mK7Z2HZ/J1cAUF+bv/i/MapJx6SHm+WtblNO81glY5FXWT96FAgDXvDmrOjAb/8u
jxv6dpwb+y52KXk2S8+brs4YLVCj6P4h+k4NeBoo+J1VhJul4mOZ7QVUhMmemRryjZtlASgFcdIy
P2o/GBHDzlktp3vehfbATJqWFNMCfYDSjuIzm6zf7mh4fQ/WnaI8xYSRdGzmGmTpuVvKnplo+SKI
oG06RX7TNxUtCNCTmFt8gocanRyXNyKpQBRMJoPbFRIop3bYfGaGpN67uIxCJL8fqWbxbSLbNzYg
vAwKfKedwk2rhzz66QA95CjVN7CJ3VRIEANIvEAh5LNOUXQQcslzP+nfh9gQMz7+kSn+c1aJRiv4
/vke8++25LOzOT1tVFea0htt9A3gNJSbXNSCor4N5VR25aH9tU1G4TI7sl/Of90LCi/h80GQbg2J
ljj2miGjiVV+8sne4/M3siTiVEVdnrdd7yCIJp5yIjX6CSyl6lLD43i/aD4Qrcxf1ZSckxI7pAB4
Q+eMNGgH4e1zu/w8ukGdGGvzw0pdfnZvJo9U5xX4Y9tRBPe4GqZdZZr4NPRSP+w+TZP7u13hwG8U
pvhMBRNlhrt3GDkr/WRV8VhR45aeHsNPiDcmky0pcReE0z1Jhr/tjaaQ71pfaMFdKVXxgLaUsx9r
6eZUxMsWZM7lfKJZ1v4vw7gdm09wS0kLUt9lWWQ0Hls6wTqb/s3hEhjmTlWJo9onqdKDGB/G+eBF
9E+5/7QVJ64AXpv3AlW65toiYzV94rFxiTwEQJ83+lI+z97FQ7hx2cosQi1cdKUwQ5Av5wObEoLt
MWTmpeo+K/oaFl5pQNogPWoZHYKvlPP14++PeL/wy76JLRd5SWnNlKwaUAnxvTDXaKTotlRM0/Tv
sMd6brqo1Kc15ZQfdVrrzXoZs+sEi0T5DvFqQeDrqDaP8m7hBUBWATwJaNQvrACxCDohgZmEiqES
SmYpuLDFr6mqGNo5g4IIewx+T+h91jeOXzYif5+D65qFrpF6mdTDXxI9j3D56ytjAQHUekyhjGWB
BuqVU86ILtqtB/tpbvbmpryutqRsni2UNE2J5gG2cafq2ks/00k5Oj+qfFvvL94SoMq6ZFdMmtli
b4CuNsHbWtkoD1WuPat8rQx2WFjZ92eD1FRvTySlFXlvabQM4O8vK8eTletjNrL2SHdwmV1oJ/6j
3ZoPsHsNgy3DVCzg4fklAq7bQUB9zKrF2mO7wkDkmkdHEomJqS11FuxvA+B4J2eZleLB3Q4VZXHB
MtFOixVShiIYYKf0sVGq5oGM+dr6s7E2p3ml/3/l9qiyHRNH4TCga4Oes2D9/3oNlAFPUzTwbxlu
0vTIgybRVeqmgSQHMVzgmadyWMDV+Zl9Wsf9Sqhx3UJJqY4lwCu+/vY/S5WEQRN3NQn156iw4fl+
oX5hRLwM1b1M41IHYg/Hl0UL9fOHjYzc863pNL7gxtF5blWO20j5yObVqtOtluwnS7qW/7Mcp/fs
YhgoAqEekoJH/m9qxXgAYlLwKT0RMKMXnfQ7oWVtRXVfeAcWvWyx3zIuMo4On0N6jDv+WnDY/vRU
9xbSyHGoIHwYDkoknXOV3FAZrPUXzvS9/DuRIRer5CgaCSHfXAmG/P38BGRLTAs1YpAHpnmQZcF6
+M/QzrL7/B9dS08vj4LOcaWfzqPbSt1R98iU6agg6m9RsVX0ywnd1QTDWqwjYxLpbc4p3YNQ8xs8
RhGBTdcbp2Qa8pJOBJ4WRN3yJVJR1a85NaJrD0M23IsakX6p1Rva6bpgfVpJTr4axlI/O7ETuWYU
86j7LSz1GTLefkTOhnmczhwh9qTjpfpXBnda/bZ7ENWEnit3BTSxLNm8hSpapcZaxbAanY9aQaFV
r5Fi2k8UNhO7NXdil2AuhAlGCozCdYjDWx4YQ1lkhyWVeASJRJyTV5mCFmSjbqdvfjG/TzD00VRg
Zupbf/JHGJtrbLgG+bouD9XgPcdbYxkEbc2O9Y3TMOSD4p8lZKqOMnxxHJtmvCG0MPZG8FuWuxv5
yUa3Dp8J+jvUdfZf6CZs7Wu40Wol9hX1bsW7QAR5lObX2rBM/9lioS9iGmTalHIfzdQ0+xJMNHop
gwwZCXTjWeHa4bGCAAfKN4Lvc7QzXI/aHJQADjnRZmuoIZN22ZV397GDORkHH1dpCFa1MHu6XxGf
tk4skMJk13iUEfi3qm/DcnuS7/d+rLEqE18QgcU0BnJ/fNtEja1qYICsnCiQ0Owc+liawT9sFNo2
M0Tb8iIRwmvwF+lRgECJ0p0a5NVBEO85zZ22jP0A1BDm9YlKpRwd8W6LkE3+l5a87IxmTjSehly0
FYnGAIsEo83PfqseJxbBITehxF4lhLXBI8E6ybOG1uyb4IdTouvQFrw360hfoJQQAUDxSEXT03y4
nFD2jaAHPYFmWwdWt/zx6RpCdijrrTZNp1hUx7foCin5b4B7aPwrcwiPbUckTta1VORqRxAzd/1h
fciQV5QRxLD47gpt9cZKM14Qlxo6Pl/SJv722JobU6dkaAztbzg8chjuFzxSy4xS6TqsDeNQbSCo
9FsDDDh9jLwevPON1zlmFH2dekCAryo/vvMGxFH/M/HrV5k7s2+U2Dxc8yhXEYoCkX8jNnavSbSL
WcH+aBwb4YjJEfrFUsw6QpjhZ0mds+9MWzk38pGansehUg3nNBC3qxQT2tqnZ8kk6NdrBcBUHQYT
n63/7wJX8iDzrRRDmfCNYGH0+FN8XnSR9bfgenOSLwJtSZe/QszViavPzap3armxY96x+jUVNw1A
vIzpt69CBUVHNoHUTVbrlq/7xkRBTCM0CawVdkO2mBV1ZjBFgRFDeoB4ZhoE3Muns0v4eYkuE8Fs
u+NVnrnhnT2b8dXqRsS+eu5Q3oGxnLGKf2hyxIktdfLRA3GUshqpQ3jJx6kXELs8vTp2sxSihFqS
RkX5qBRQYUEG7oUWlHLu3kY6Cq2eCD2YALoqDIgfCuUSAcsDGh5p3wjrseDp7bEphQEIn47h8iaC
zZr5fPs6rri+vfoyAa/m0bPbg3pWXQJ8GHb74BZ2Bl1jF18mZL9Xf9dkiNiS/eJoRs3BtvL2rOWL
xyb8Rl2xaNT2FqEQdmJ4cwf7UlveG3MjViKWwigu4DRwOk97hdU/dJEOjxo5UoCOvqZxv5vS35al
k7pZFWqeniSUyekmKvXG1HZ3g2ENL8xTSDHuj+HcwjdXoVEe0KFpi1Tb03KBr5tGntU/8D+D96eE
f16a9cyWk+56VRRLD07nHbc8VD1ozCX4/XxsaaTXTtBpJSIeOmP/kfVvfgCFOkZQhekQDkDufKmE
xXlNoTU3eRzVwIBzMoegT2cDUJ2RP5JRWuuqWVO4rHcT6TEEHoW2hFz54OIF8FHJJBA3Ro2XcYBW
5x0/zu9aUDs+Q3cEWHdzppayWF7MhitTfTxBjgUv0GlVHeWW9e/CFMIVgyzOiCp3ZnkkrAbbwsbE
euUV1Rwh3X0bJtMMAf6AcTmGORXfDWNV8n6EnI6cKvgEqL9TY+I1Mk6MmUL5xKzqUCRa+YDiXnOf
f+mMkmKUHrMYfM/7y22cBxdX5igxpdS0Q3z6/nnaaueKWgJWZXsbpSa3Ej5R7XkhiU1sXN27Yq9R
68qEAIzwLt1RHmDPJYnzazk4Q1ZO5XApZ/v1FPlQRnCiA6+kDbEPQGQhKLGxp55iYcH1+HmtEasE
RmeBi1QpxITPVGwm1V7jGQY/7mh+jWW3Spdx/Ovhp4sLwuD8BKHo4YyGMPgGHY2kYXS9jMMqam4Q
BsnZDe3KV1DS0wdNa2zyd2mvL0RCyVa/F4KDJ8Kqkfj/Dsgp9ApV0HCr9DAi0mfNpQA1cOvhjGq/
XB8ensufQYIxfbBNJbfgDztG7n8F1L0MYrb94TvNSxo8yeDvLm7MOkgsxhRyrfwnoLvLLq2aIwMQ
cdPtweLhQ5LwK8jB6S6iLnRIJiqhgQ4MU+pnd9OC2Vk0Qz9mv98XPyBMZ7Pae81SrvOJ8SQoMcUC
vBtJij/sQpRk22mh0xCNpXnMZUZjRFtid6bq5rt+P2U48a1g8YeIiLJxGUje+cZXVmFXTUDcfno+
acDai7dKO7vas93ARQAzTL3zS4l0F48ddFAple6N4eZwghHJvXs6ac0zhJG6QtCVHTnY6T7Ql+ap
2iz3Obsu7X73S3f+j/FGKt4SNFAojWDQdaFfg+f2sqNjq1OymblHoEPvs4+sK0JRejOm0zazEDqp
cLfMTChBaMNuhh5T9fHa2fmtkJgzcQVenHt+WoBEqHU+lHOj7wIMSEKqqSj7hjNZgPBkOTGBD6b7
1YOaVxDe78xUpZgY48PedqEiWKSofk22pi+pEbI6+OhYlxIWViK/ONsrwoUD3E3HYmMDEttKiXuH
pb0cDI0hXfi1qz+QYfxOSg3TlCiF/M/fVwoYsl8E8OAkCn/xck8jAE6dsSG233kr1g2U0j7b1SSY
BFhqwr7RmwQqDU3BXhDpFttGP6A8mcrIgkmEEFSw+PbrUEbAo6kaLBxekYuoEaNXnVsIR8MAB0pD
dBxReFAuzraL82GulSq3vrkhVikMvfm5qxWkZH4CJOyv7UUA7soeKduoW3Xc3gY9ouKVvUBwz8+l
GYzaWT57udA8RvYJFLMT/iUDKt+x4OU/cci0P0bjPfaCOQTD8sGJqdvH3TMqkDuyKo4r4HxDO23v
/2lK2PUcAquWdLW0t+f6KC6ecQwaPR/tMS/QT7QSsdCcczBlRGPfz0vZTxA+SUWkz59vG3nCq6xD
w7U5BuAY4xpyKMMWv1E6fK2Ov03s8kCY/4PyZ2z1al/oOBuDvItEgNUPb44j1zOADFTi+/0aLMv7
KkAzKUIN5HC/VA/V/0gn+lz+k1pOajzRrLnZZg5+U4jGtaue7+mM2grfA9tu7r70GI79jzc4E+2m
Q64vMUMQMNXgb61YPwXQfglHWIFj/QTbQjPDO/QczsJc6D/B5MH23Z122dk59aSIh8eQApOVNQpf
GKcAm0Yn5m9fa2I9KnwrspvihrsfbZx9cBr2jQ4+/Pqy6m/w4rlvPqscs4DKcPMp6eJj8ut6F8E/
61ziETWfMRzJCOd8XcCHLYWjPC3jMNKOe11RiZ0u6qQQr7xOonYvbbfxljKoX9C7UcrYOx7Doq55
C8KxGupMIBAK6ywq4Wb4VsnBXTJasvSRs3psR8WEASqbAs0rOEbUJHBIs87LjCXmguBrtrB/OcGG
oK0+JeLxYONkmPZdrbK4IuR+k7qO0W8sbwYNgfiFy0QzMcaEl5KYOrwTJmyM7Sz84IUiWFeLDHl+
3PyoP1Sy/trnYxLR71VCIKyVkT6OTrgUwIn26W5hrFm8fg7NpP3wgiaHP9q+89eAHuUSuYlEJnRq
Qm6Yd0/8OlwEwCeqAXlaKeA6upEWRohornDjQ32Az1Mup1sxV0bdj6RVbslViXaRBxv+qFkE/MQd
+MlN9Izp1uRzGR35p2MDkZU4BQjse18RMCapYBwc6TKUfNko9IOtp8a6o/rjuntmjB0DqQzpNjXU
U164byIUefag/dFcS+EQ2km6i2nk6IE3QbeP+nTaGGI1mtIg7lIfkEIpes8wMvHAM37UFzpsTd71
KviUIRe92SnqU4xjiQEffFs4gf4nCR7glNLUOELqXm8dKQ0IyVhLnokU31y6sRtPue4c37yn1vXd
0Hl4QVhZXYpjL4hz2aMzrrhHt/mSJ3mZADoPSW5bqTc62ze71VjUJjOi8Aasa779vJaseCgJYnk/
ul23aNBongtjjwclDIaUw8tMgDS5a+DrVemEvPGz2JPpUdVy7Xozdc3tL7LiNoPdH5ujSgw2l3fa
NdmZfKywpuD3AFyFqnD8mgGTWAxwgfE3b5/XXvoMNrEHFyHutDXuWUptONyY0L0eKbGUFax/+4gD
0PaE8EM57gva7OItg4hZt6WKiYZv/AM9JotrE2YTs4e1GSjEdMNBJ/UA5i0k8uURtk/EpIIBfFcm
oSp05sE9ctbxuOISKOQQwLVWSwa9G0mZWSADbJW7US0YEGSfADHd1nmcucW/VK2H/Ec0AL/DB/Q0
bsc7LlxDQqNRgnrTZOA6WC+DZiu2krzpbKla5JZ4fYk+NSmqqF6cNdb7nZG8t5/BJzO+Vpd0Zp/H
ugaNWDpselWn3kcETPxf4kc6/98w/leaMGpPH1wIJZu4Cfls529eQj46FK6Vm206okiCgzWbo5Aa
elXIxQTeQUHpQcgsScrGFFAQR4Wt3Z8XfxZeilNOrJndOYTJ4swf6n0DZh9Ufmm33Y33BugdU01Y
EF7s6GcJi0iqEFIpqNgafn2M78HgKi7+BNXE3qs1/Lxkmdn6bpzHQukpME/GPqjr5x9t+0v0AiqN
FHJM6WDFfiU7KT25KejmIwocETykcyLWlnigZSSLuwRVAp0S/QnZRVbuQCGGf0xkhP5iSrUvXLuw
ldbWFsrsVwW1MDNNcpu9ev4N1Eg+y1acs/SWdycjKr72gHDvXbTywj7mG30GRpFi0Hmrqu065Njn
7GU0tsjQY8Kw0vDqCe0XL8ax3WqW62uvrwxrJ9kb6ueHzQu7qB+cstxJhmmlAlbHcHvohV7VYNF5
baWMEC85OsFMw/UE9N4kQ8esJYatFrFF6RRpbByEHxuh5+ZzbPTUSFTdMY6QfcTk10tYFWoITraM
/Qu/Y3b0eCeTsu+OqlZMQkMcMMq1WOr6bY4c6O0uAhIpAqdeeLElmci3ZhpiudO4txBTG8dj1YEC
h3v2vbLbpPc+T9K/PlrDQDExTGXndddgH8zjrOMMJWUWpzS9Utd8J1uDWkOmmgT5nh3ZD5rFnRy+
820Hbo0Nt/L0JCqYZeq7WQYeVPLjjopum2xwQxG39wrwCoTaY+C/uCHLrW78czv7o3m06MwzlBRJ
9f2YtWF421jHS6yBz63VGN/S+yhbyzNlTKjj5iUWqGAOJfugR3Z/HaV8FTdvSoqFKn/sQT6zIDBN
4pt/wPcW54n5iQuTTwFb8gmkFhZxlOh60H2W/2jYZsw0GRFXmagobPLhLQXaCC2z90UAHkVmsI5C
MtzUTnUp/1kYhMddEnuK42w9DP2CjGC0GGSKC4sfw5Dm7SoDvJ7LNW9wyzGkgwQ2ILijLecA3FeC
czQzwBxoW0s9hU47hLekwXfMyQymwVVun13h5hboatiP8++mimhPl3D/PAvudFeT+Ce7G4xMCpwj
3EGnWVqYiELidajTTYUOuvnRD+CsS4N6v2zG6KH19i/QcyR4NRiwolL23WYcO67vaIyuzTmarBGv
2erDyCABwXceGgTCsQNKn4IPCPzMrApNriS6mE3PR20f0Fwt6UVWy364cMtg1fTk/qx/bBxiXE24
vs9StXn0cuTe4hZD0jCVeeydH24OAZa1WQ37n4c0fxUWsGCVSEx01tb0Wit+/lVRhv0klhgfdxgq
2SJSTfRBRxLR+oMh7DvrpE8pVRN+WSNnfs7hZWkhjuTOcVSRCK9WVBtAVEeysEK2cRqcKFMBkZVY
7jCjVgLr9vbBMggRAxdTKbhywkwZXvmbNwATcdag8w9uxHvFIRtGzjYUmxpS4ZnkFuMIj+3UYB7g
zlQ98Bq+5JjpXAItCwNKxVf2OrUfb1QpMk+sWNqT2TLP/xVxcruUfHKD1t5i63hlmK9UGfW6y890
d4w0ORP9k4TUCG1aWcbtB5b3BjbGhBJRWCrj/bt5xd/bsquJKDCM7H9pi4qPqT2n2Jxm+WFNV/Zn
CsKhaUwe+SWBdI5swcrM/ZHTWSTnxelrWRiU57ZGZjEtnwFBHluXD4A8nvWZZSpCnHFYwXN4TsJA
09A2eVeKJiFJlrb+j/K+Kyx5bE8sBhE6kCspIBFUOkQNCIxOcXrVUQ4s6AtJ2HN9VxbR1yxFV8Ax
+hOiOgivUqWYYr3lqODcOK0t5FPlNbqlvwFXG/5H1IGtRKJGQZQpDXlyOokp+tRLJbz8lxflm6NQ
lYcz5dx0uTP5BSM3r1CdqbuJNcCk/cfIqvFaNADsvLmkFKcd27nUeopfNledKb/y10IV4Yd//bdI
bTq7TbcvosOV2G9c+5AJ48sG9E+H/iU7wxF+99f2FEoNYFYgbKP4qy6DAigPn93I0NWURpx3z+ie
PP/+GogMvFdyEAE6USoB12ByQYTyU2LybnebX7bsCsybnasUoi9lrz8Es5qG/3aABffBEKn3lMCl
X3jQ5N5RroDhDQCQ/wKkRCJnFBk33r3vUKJqMpX5rEeuv723sbStC+DQi7fFPNrK0FDyXOE01e0Q
TE8gfsOI+wvSHF8z/Otn/0ajReQoxDXANr25cmlQDMl2iKD7SsjLi8VQryM4gRvBz938U/FinUSG
wUSRQRL2//k76/8GVASJOHdhCyT11e7vlkHn/1ZvrI77bN02pj5f7sdktk27oGPVMxeLRdWELRu9
ujlegqm8D3E9vRXxua30yl5tl5AmMAxQU4egHFs3+wIMzoxR3QBN+KEfSz592KL06p5zWkF9vXI9
wf+Fbm0ecQMVqdmajxuMiqzznmH1B5GcrjclrYYBCi/Rynqf+2uHqfwAmeBLlz0WDhKlF6FMv7ZS
X9bsysfdwZ5G+l8wf8F+fsRAtKn+8XhRTbfd91NUES+7h/B9phB00ohqVjXHjv0JdJNdAVvXYogO
ofThqWOnGpxfZ3mWgWPAEs2Zlj8MyS/IJ9Z6CIRY1Rs6ygvPUJO9QcXJtHjbhg0SKvY69y2kll2g
wKF1GuNaOZXnr+WVL9kaA1dZP/Sqn+thVjNBEeNbuVs3yBob4nDlhHgo05mLoXlX3CjsqxW4k13B
lM26N6kP2Blne6i4FTVJ0jEwtdn60+HAjlFcABfg+A0OTLPgJv/Ccgg0q7A7c5ghBBuiM1HqQR35
e3tGCz1yPYktvIfqLYL6IRCGJRBP36uyLY0BMu9tStjioHosWTZ0WIT7SfxGF9Nwjy1OCY6Q+Kia
J4l0MQaYNhTSrAcf8o2TcQgormR+c4bOsZ3iRisIIMoteI8zrjbT6coQOxN9u7JqtavSmVQExUsO
8bgcToPCe9GPbXIMBZaaEJazxSbyDB+oWRXYu0aUxZj0e4gtHRAgeoGOxCUyXxQaFnd+tuyLj//7
CwOoCQkAIBGX0dLb7oGe2jeJ1tk3iGMuab16yTTU3IJVa1Yt/DQo1uAMrih/vsq0b1O1JKathApq
ux71h1ZQfOpq+dSaW5I/+NDmoEIkTjlBS2G7HftXPQdI795PQVjnRoFn/BXhIqsHKgE7yqIcV53N
yHb6deEBHA7v2s+XjEs3ueIpf+bqx9+jLP/mp/6gEGIZbSNjz14wfATZSP6El1COJ5WrqA4lI0E3
4CI/I0an6Vfz3vZY5Lw9HqUlnzUg+Stl/RMekoGRkwa8s9LGtffIHpbTmliVHD1KHcoTVN2ntVsV
Ze9Dj+6uE1csC2sq5b59KQYpGb1j7/4p+vm8fIq3weIMppar8YZeP0+HuUB00aAh9wyv0bNVZCIU
hoZuoICiqQrCVrA1m8EhQMoBzIL+tjBw9Y8uu8DOcrWyxnaTUOGFdWmWi1gvgnWg6S1XQDstUiTx
6fnGQWg1XAcgZXEIVwdJvFJSD9qT46A0N9QlR/RU19zX/if2Y4l6wmhdF9LOjkkSM0QO44j/Y4AP
CZtTMQ5Ncjg7XeX33nen9UmqcYRNcTG/v/abGgpWYc0SHm3LxyLJTtmDET+qmT/qDZi4+lisuYEv
THe/67ra2s3dX5RufnbCYEzADS6mK0736qe03iFiUSRboCBCWSpd5KH3ygCtMFPTrFawMi9/gj0Q
l6NL45/wKRg9HnfE8SdJYrJ8zKZRp/e6x4lE/XdAWYcNiw97+gCmUuj9HnkX9+9JKmzBFjwsB0hc
2DAz8AB8MaAez59aI80goO2ioW21P+Uku1itiIslmImhwTq7brV9FLsgVGqcZ/OJ3HG2oYRFCDHs
YxtaoBzA7wf8OhvxF2BscZXXC6RSzym751tQev/X7SzJc5OxvQs0Nwlr3HOftMOX80E7gb8y1v7T
BxG8woq0HimqtWduF+W9bB6C4fugQ2w+Z1SYKzwO6m6/HuH/ElCgWy+b7/EJhTuk8XEIgGXnMgaW
s6yAtZdQsszmyYo7xCoswPwbZKZlrbMEmoccA8yZXd+pGFzl9CAlUNCgqu57csffXWb8A3BSMWIW
IX1SHBnGp7N2dqgAwDgd1DCzvayKANrUuX80x8KCuOXbAFwVcH2ADFjaXvoLBBzPqiD18hhErC7C
AcPyNu3M/P2xnoUKqXc/Nnz6e9pzTopvCx/Y+0wD8P5toJVHu8P5M0BQsKB4Fh1VzUPE/4IQ5h0N
rBy4m4teAJnZI9IwP4D6TYg4+u8VjOyVNYi1Q3OFsLX8w6sIN9TlRTU6FWUlsKChSbF+T/WqNmI9
N0mHvyS7gMCa/UlQh+SJnhVUWDfAoxP4CIZeBS0sEOUJHQL+7YBhqdUvbL+es2xoDlFBBqogyxHu
aeFsCSj+X7foN2xdI2F9TN1B62r+kByxa3160cGfBk/4Utjn/LHO0+RCsqTaMjTzjWp5xLmIimxn
doOmycYd88k87WwCQ1UlYH++vXYJs1s0hbDoo/d3qEXU6vkVbYh8x6mNDzPWsWC96VFwMTCbfNBl
+XzeU2svfouCPLGXe7hkDxKhqbmAXKSkhbKdRae2h7vwVXGpfHIu8FuwqkNgaIMuFiT4GzvKgS4B
97WvCM5ouyWq4r/GntqzXH8gb0VE6/hFfUbdxMTdH1eIIWhObLrDqFv9jw8cGylZGwN0ZkWPeHXS
xX+XlZCibQZPTpFUxk2iImUFSgwi37NSDqzpd+A8LoMb0tvliBoXVg2Cw6G8wcF9RCCV8g2a4Ryu
o+uU5HfpU9fUDBNfWo9WTiyfOzYFhsk+BwLIO4lWy9zOhEvii7fRjTCTzMZM1vKTUmmQ8QGLchtX
gp2CatjoPJMEgRcwIM4BycMVPHnD7jOUbOWfZK2Emx7rdz7Emjs1j1MvC/Re0/IXvsTgP3lyqZ9j
OLK8qynkrcYI5mlZudXbPkivNXWQA9lT3IYQg5pbjDCjofTAjCoGRUyzHU9Zzxps0zWnS/vRqEyJ
776a4nQpt3ovbtC4FGwPYs0TVQjM6s/yrwmMJ/pha6bxZFzgdNtGUap0uRIPSWUewUkO5Y2s2ySb
6/T3vXDmtC+DzlrAhlLlTpo6v6ewpU+JJDhe2SjXNzVx2Cxk7BKQBh/ztDizcksImSXlPdi4vzm4
bPOXyWGU+rauU//uneKP0wKptmHFtjMyx5DVbpRWnBX4j/BP+D9B/4ng+dmg1ZLqTHv+zqLxlqTb
OSzmnmTimmiGNqw9hYW/IhLGEWi2cZSq2XTom69FmG5REh7EUuogHGE15203KsBfFz0nBZkz2oVG
uXh5gHJBrOV9EWsOKtCdmLEjbdMzWIf8LZKd/tnWAUkx0q3HtSE1By4rweOVn6jRDmihE/pqjEOM
YJZKusA6jnqcG6dfCdQdq5gCTNwHT+wZJ6jFlLj9jutQP9vO0/sbaiFXbQcRECMXIkrFPaS+LFI+
muniiYuVtYVfErmw5hZp7RDBTMzL3JDUcphXukrhzE6zV4z/GufbxTGJ+Cy2wZqMjRSDO4/znapf
CDHq/iFlESWOdSGo2rcjEuTlt448cvTc0P/UiBzTsV7w7ChPwyB3DfsIgD7tijwIHcfEA0bafiVF
GFRl1BjsHIN7iwGwGgz8oWEcGe6wP8BXAG/Eob4kzYkDpBzGupq+fMUX093XCa/L5hW6zm63e/y0
vb2LWBzkXPyrhGjT6SJSD3XX00/ErtqEuogBLMuuYAfkDBgO2/+qUh+dps86M2pRljsi8d7r9IKp
6MQiP0zTwVKk+FLo0f8rXdPCp3TfrinFxIKhCSoJAp7J/rQ9qeLilFZR/xW2ACQJ2isYrGfRIaZz
gZxreyAkqnP/R+h2MLY8Dv3RaeJk8qY+g0nSaQH2BrA86cQYh59ZRb9YD2jxVBN1i1pe98jwRKDZ
5Si8pNYwuy4PtYdtSb482WTcgR5UbhVwHiPGBkC+aanpkicwK2D/56LkCuCQvrWw6xZ+D+fOot/M
2afsOvvINUEN6Aom3sRQjDmVApX8CIuFn+zuplqxfcP2MxK8pDu8osjKhhPtn99XnlzqmIa8icqd
WcvUM1dqZCXDDcic/7gc3T8gGvi43aUZCM0f0A6rfOu3tw965ltrs5/eUTVGxVPZjdEDeDxFv5/g
CSOtvT2aiQbJ/3hOhHHDSE0AULJSIToC087z70C1KQCR7kZdgMjx8r9eJarbpVvefMwUNQnmgJr9
/QWOmC0amtaUxZJSZiX5qqJHmikP6RNvQD1jyPpxp7LMbg/EqS52jvGC7aUsD8tGSv3q0iMC0xke
i/rXpLkulX/bGgQgko5BONsNl6nhpXkCt6QSbjes0+OlS1B2FrqpLXw0M6J39+yIbt1bmTCkb98J
OS6Ck8jlZeS1NzKfd59YIhgBmlpSJRhG0zaEwlI3SAh2rpRsIL/Z22iKSFvvnjRSutR+KO2/vGdn
zWR1UPsl/4kwoSHHOisDkcdQNONvwghpkdpILWH/MybjjaR4EGOR481qCd5DnqcWedaEKbwBIPKs
8f7scZkDR5PBR/il98a3bdy+zXAV0q2e4EyqfFtKgIGbeDCO0i3NWJhWCyi2FPEWS+bOVaiyYL+o
I9NdSsIJug09b4raAGT4/OVHlGHSwvJs/5x1PlwFawlyQTTVmtGhDNQd0yM6meAsumYQi/3m9z46
k8vejylIhLVRkmztw2jD8YUbNP4t5XDUotT9lckqM7nYPkRss1myfBnphg8gQO9DicLyG4f+ULBl
9wRm/7c6IV6Rg6rmD7H8D8qhxQ6OCDrV0w5hElr7tBT/jvts9cjFxgUeGDg212PK6IwGZCBQo1iR
NkXrQ9MfP0zf1rcy4+dZvq8OL0v5QRiKQ56QFCvcA2+05f4hkLD6xo7B0TlcI8kjTJTUV18zdN2z
1mYJcWNUtjYQlfvvT97kCnf0b64nj/9XtvtPQ1D8gkz4ebi7m4ZlBuiYfnmeN7wJL4M9VUGJGi/7
Ef0SFq4Yx/+iDSoc4zkACAAewtdwt20WDH8cw2nyOswHwkzAHlcajAWPUtJdmmDMhnl3VDEbubsf
63GlBAPUof7DBGoug/0fbgEICAbmW6OP8aLOMYr3xXXrB78a5XKm4i1m8pNQCqoJeu8T0r0LSrR9
rukZ6mobgDzmq7e/vNynhAmjumCYn4afWvYllFEjeoGMm1eh5drB6gtZhlpKXOcB/k//n2IEeSVg
mu3Kqiu5vbckYjfDME5G/r5lKuMkD9qirwSm42eHJ2TogSK/6OHP4zxrBP4ZFyQ0jHiLHrIulCEP
ftjuKom2OKuv06i1IPi5ClhysTYD7Vpz2QkosTjMzgYw4sH5fkQKseqihhHolVaGKfqxtSbKCRud
zWBV/yRBB+7hh0FvnQTyLEe9qU07N9X77C7KwPkb99rFkJvOXRY34wX454hPRhbAaG3PXKIe4j2e
mbkdxBxY/HwqN+iM7T5EuHKkU/sfeyln4WFq/XoH18Y1yC/anD7WvjdNom22BfEDVYrxbeHOPcbJ
+erKxlsrYza9MUxQoTHMVdM2BRx4LU3XHi1z6sF4hvoPsZWDv+B/csfzhMs+72JOokxVtTE7H4An
qG4/re8YndwDp3/WG0IxlOXvMP6OIbERTjgAv431Z/+0WLS8x+BefDGpIN70RgwsfiSomz/yUV24
IOK4zrEKEHfKMCeLikE6kIZWq0QhIwErkdmgOzQUGPQMGolTYZGPTZmvuYCKBqvbV+kFoebMEUrW
4+sdzRt2nVzfNCZg+IXWR8C826rykGu1mAsZTCrm0/7uMhjuD5fl5Xdf/rGUOIs8Ha4cYnQ2fKJn
Tvphtk2fUZ3plIO+TAEXNlVEqQZFZ2PHspfk4LXmrxVyIHVFhRf6Ky9pxEFzw6dXY8HsiFs+SCLu
UN6FZFG7VG9C6DEpmyZ+exwwfALZMc84PKw/ru/Z9Wy13gJr9DjRZWrpLLQMvO0GC81jfsTGlMuu
44pkILIfMwBR24GB9uKyIUi8DbYwdPd68KRjfwvDD2F0EaXfZd6+h+GudPt2p5o3pDNEGaJR18Mf
kEwnVhVWWCF/YjEQX6Ia+v79nccesZTluQCd9V2dCY94vpvZ6EfMvRBagqGyYHpp18rHrbpiMsxA
i3Y+fKsMVcnFwfJ0hlVHeJlCp8xN2ZASVbSXCrfd97ZR7rlC81c28afCZBstiAe+BUBs1dps4Cpq
wMZOjggHJOG+t+pakDoiY6rrdpeJALaDZYFw8km/pOTHgCQC/7yRmiLnlkqI8W454zbxxKIhSot7
Np4u17aNRlg5QGCzCGhuJ6m0sxBQpwvUlM/5C/Hs4+/XPw17tyK7vGnN8AJzVEIn6+AyGNAgOuyV
J4DDPJF/hWYitojHdYMK3X70BLvrQX64oKkjrpvPdsCmHN/Mg5h6jBiqxdcLtkpjW5gTrRZTGWZY
vFSe4h7f4ydvenEPhGA9okrV+hZ7DsEVRh6BQgDr95gkZhp4wgKZHqm6wl9utCZlze6pWH7QgcOu
gwRUjBJEtwEmMqgl0So/VPzNolCDZ4vKmWd4I1vSyjcUOE8DNtLvTmqwetqkmSUV/nHC8BMGrJm2
FpgGPMIgSdmsCJCNGBZwPOXDHH6QR+nzgmDJyNXAuJ0Ia/4ES1otJdEmb8TrfIu1ZWa8cU1vsEwy
UOucBPDS/cgl7Ao4rLdbQUqCg1EDP84+kUVBeH1Hw56VnlJn497iE8xpQk+GysMR51YSBsElhXkx
ivUlhn7STYEXTBqhRf9CIVwmOCQdOkuruH/4DhIXL4qaxQ530uTCO9VOfZejOehjKwve2bFdE7XL
cXj0FK4ieef0Gf0/SzcqMROwVwVaTZSF/sHCzp5hyoql1OD/psTVhqTZciaHS7BOUye3GlPRRzIM
qno9DNw46vwwIb+zUTS4ttVGYc/VAZo5FkQiG7mQP/6f59sF21UQXpI9oiKM6JJO0fBVIawvoudv
0yvAChr6imAmLksPHUUizTiZKVWe++GZwiWVhgKZiRERCKnB6F8XplGBmkFkPvZB9eN5EFza7q9L
RCtnjkk9ZECKSWzZ+KpzkYIecwvsv80xtxlPMqQOannxZr3CObS252kWcEO3zY0wzNN5pXt7UvcQ
rDYUoDrE2Kp7e14Ywpi1DgP+blgMnUs0IkXH9zHJXe/zLufY5h6bz9aB6FUZTC2aBgoV+EX6vwwu
KgBYwylaMSFqxMk3hrmUSYl5n1Ued1bR1GIlKvTj3o0ZwQAt2LpMb23+SWjEIBCnWKFncjmQaqMN
uAWNib2RxW7jmd0TbR+BZprL8zMoxU5ARgTUzhT0BLbuv9GjK83d70rsc9jjmwuEoyuQijs1b1hN
aon2FhBuQuV59OhuAGRj7JMHogZ5icQvrWHsxbNxId30vpEHQDfi4DqkxIue/sD+Ehvfig8YYg9Z
urOGcASCaExoaZlcaU04VHuMWBGh6IJwkaFxE+fg9ZT8s6NIaYBD7bYRvntHahPMc3hevao3y8h6
Rr5M/3DYVifnfuFwBOnhIkMZ9c0dSbopznY/VztGIheAKvfeojUeyprIic1DCjgatAE/lqeTTaWu
4ovIqoYEc0Fu6upAJZjpJz4d/wOBZupF/imI+rOuJvtrAy7OzBL2nBVD4iZ2h9I7q9ivlMV38ZxK
pK4nst8fcdRYXiI+sQnuBG55aBD/MOgtWLTT9dnjsKonHcvO3u13ihSLQIqjcnY7R6dGWl4jXo2B
e6qtTbjOFCoJVFRXS96YeKPEMc5l3x1KqcFPIKm8jHLqvuXfz6TnVcGPjHWFiDxDu+DaDybZdRuL
X6i07Mf/uYdLxj9ExjexoE/wsaxnccijonB2lP384LgLVWtuOjssFYB6QNRhNjO+eF8p/M2hDoSB
V00d/9idKW/Q6UchbkzF/B1xn61k4rEWbLTGaoRiN/eUHmq1SH2cYUVbA7iid1G+E8GO09aqLcBU
a1Tk4UMm/NZPR07T4Mwol3flNxmqf7yL9UwfCZI+BSmPhZ/WN4OaG8RL/HcXSvbzisNiggUvwgZ1
PO2QG6/nOwRCqeQ/UfrWP9/U2+p/z6t2SVgLkUw/i7ZxE6WzNF4rC8PCzgbEjXrad+SfWRB+t/Z+
h1zt9f8NYRKkxjXwraDHxXzS+pkqNojRywRYpSCQuZhcAiP5v41x8+btoHANykT9DyObVCs2aNoJ
eiclNahPtM6B2lpLy0emtK4UPKodgJf3zd4DQp2JxJvOKr1N81/RJg6BP2URD0DgrIHEenE4Chbo
OnUi/A/mSIoLJKX603vmn75gVmkwGlqEmUdmKyMUc3ky5gBWBscdIQ5L9B9lNcuL80+AHeYrPAjD
7dghSypZV9oZ2VtSm8UizSJ2F+Pl9PniWwXo9x6WWtZyvqUt6nWmEjA31UPp18DoX4CbIeQbmaCj
lXaspTBRq7Ts0EuJKn/q3BlEsAu4bL3wYCLORue4+p73UxU2ON0gIiGlgd81+e8PmeI5/4TnQQt0
criwa45fthq4U94q5bye0GLmzit30bEClOmfnkhqy+aPT3VV5ApGIBCmepZdFJdwKgWI9DhQzboj
rxaUfDuLTv6nXTj2pkd/QyXkdCC8/KrSAGTic4opoRzTJMLciQefe68TpE1xD5y9WUAFupWvaoGW
ePe9Qc5Xa/69NkAh6mY1XpsPiyD8R31RwMgR6HdZ0c0VWpgJl6pjhh9SZKwRW9Y8OCtoCKvByXi0
3YAPnppIoynS2Oy2a45nbNEjn3kW/VftN8ytoWBN94Se/M5v0+XFYAQw+WtpTChyK+TxhP0zXidE
WI+BPswhywTxPbUBKwdapCwNKLKpSyg0zfaEubgdxYHivdKbb8iINVzQN0Ebi85taiRcd4C4tigm
G0pKyry3IziCT4+JNkbL5qHPW+sGnVeG/8MGaEptRsNg7GOdOmtJaIm1qs1tQKRA8ej1fouAJ6Ds
YUoDFMU77x1AxQAsLVveNYNJL7qXQyZgZwUTyOvFQorKXKGQs8iRQFErJJHrys612j3guEMh26jb
ustFUQPxvzDh4JS4a4RnnRDGk7V1JhL00GhUugKHBvn4WnV4DCP2u4/sRrwRIP9hx+I6zzrSZ0Xk
D/Pn7+QHk3S10eObGhzo7rCO2sZCGIHUGiP3XcNNZwF37KiGf2PEdDpnHV1Xvy2oehPAcNodDOwP
x9Dji65NzfjoGAJLb+MBFwXxABNsJ0gOhGODLI7djra/Us33TwbuVP5HwteA3Q4rK+TztMkOHt2Q
uOgpLhaiXexnHUJ0dsPlh2qhnA+BqeOuBlotur/OiM0VNaR55KsQdyqQwwStM7mDwkIsys3hNE8b
GUqEUXp1qy3UFgf1he7zIcrtzr9RPX6xxRFFpb5FjMSj6Yf4aL6mx2cwBxmORQZwXNYyvA0xQ1zo
xuXY4AG/ve8pjf1d5EwyR1CBpCJwDF2+1U5k0HMmAbFFNE3rF6tFgtiE5Y2rLaoPWm9OZtS2T4sG
xOedY09uN/JAYveakLRXRvlZESSCzrCI3uhYp6ZvChRGi9oEC4qLegCqJ5FHlsCSsaBn5oZVfZjT
YjF07IL/cbnW1gY9ftKKt11Gm3B7GomBYqpip1miec9ti1lhKySKT7IpxHjk7N+hJzwgApFpkzr7
7jd5h7VvaR5tcrAdWQFN2nLAtO1mqmQ7rOf8qpzA5ymSlgMAgkDBSK1GQbNzeu2fW6Q3AEVMVuCU
e90DD+BQQOlfBWXbNmV/513y/Q3nxCg2EamquWQXk3aqLHEYNw0eKgykoO7/48RGQlz/PsZYK6t9
PFm/NjZhw1wq67H9Md1Fi4sk6t4D2ZTsDnDPJVnJqHE8TSuMBahDCUiyiivDXcQPGwQadnT7T2rH
YAx91EAjJgcKN9X6wQCvCFUlULmqn96Q5k4Ron2+iIWKtIo1zhp2Xd893QrUUQC6dueFt3xcTMi/
8ZvZNFo91FMs+TQ682p6PA+4nTLMrFmL5XD3J78MmIt9aO0La0xG0iUlfQtw1mt5oz8POLvbWfmU
egjuHBGEeCA0DJN664XC7BIeoMmEiTAW1BbULp4aWUJID9G7NAPWOo0d2zbmmp6Hcot6MWwT3/Q6
6kiTZK1nF9T9K7IeNF/huOeiHiKJ3sA37+b4zJb7Yy/66OU4JxQAJRMoPkIPO2sBkoqskMtV6J2r
nKE1D0N+QKki5UGKe6HBgXjPsHL/tGJpUPaBxNGJy45dtnGCfjzcKB0X5I+DEiPfpv6kbOKjb7kv
UNTgmsXke0nsTshaaiZF83C0hWtg+06CaSXr7vsv5p2XDyq0cctXf5kJfI9ytxrDfT1+W3HfqXrM
+Pm9AAkj6SZUfYOx5uXTDJZKx9aoipLnYerM8q2znRkgYn5rTAs/ZO2UrGvwKQckPGAQnFeeH8nA
TvTEo3vUQIwpSdblFe7khvyxdWFCDXSrR72UHB/idnw0dPB2ezWad/IAclp/30lBvFID2Q0wF33w
akSQQ8FEZfRT1r17Yz4T2gDfEofDoyK4zD5qPye6x0I9nZOqMQTc5iY+bK6Ku0lA3/XdKEwgN/8a
EkD+Wk4zAfJJo4+/8WCSxeAOd35NizDSG9MU0dWcw2N9ud1lfU8q/u5j33FPUMYW5x6+ByP2lwlI
bR+oGO4iKtoS9I/aXGqVOO772XZGRObQHvUJU4T5dm6qKV+pSsdFbG6MjgxLWsNv/LPbEtZTQJtL
ICG7wy6cY/ALhsoTjyK/j8xdvhWD4ZDw0826jn/RE2dFcKOpY0jIA+RY4L8k0/C6nUgCd6+scKLm
+buQbzRZf60x+PJNZMUF2id9gbDO+PfC+NAGVNrn1cLP/RZc26kX6BrYNd0mWlI3E7WMXqJhm+I4
vnzEORn/G2USdGqqg5WZ9L9fMa3l2iHe+a18ypIyE+YY10mER46dAkkdr93N08API12lqwoXiAsO
R//XfGvEuZr4rL2jj8MDcFQFvukvgLCZUlmz/T6ALESGHwfy1Lk8NadIPSHPfdnSr3P//rQnxlIw
kmwOcarKx6A/AEGYiWOEG/nDwRkNvNWTpr/Zj21Gls1TWD22KNFoOQGhfWlIE3DkBKPXaES38vqP
9d5uIHEs2hi360tU9XJsyFLFOdrP8bSFtkVht/R+WcsdW2urbbrNvyEWDOvoekD4FmOLuPXVByuc
qYAYDaLr/6nViPl/gnbNtXFFe3vBXw5wQ/AQTzgb4t3CkdF+Pyj8cCg/Sz7DJ3jVmM6kWqsCDWMq
X2vUZVLvtD6CF64Iiq8fLUyz1pXjuz6xok1Hv5hHfd1a1b3ZLn/P7VZ6SeiQKi+1Ov2iJ3abxPaj
GZWK5nVX6KndtnBawC7KJ+OJn7AhazmbmqUk02WaTuwJtTD8XMlEFaM90JuPZqiPxLtQBOY/JskV
k07uSv/QaFcNsI6HJzI7jA6tzEvh+JjnnDcfjokc2Ujd1PaX2dlp4CbqrS7v3fihbN1JbZ1/XYb4
M5MrefOGJkW2NDAj52h4WSBHa03u/VBAn2/JoWHstpu8DGXeMnTXSZqUr6nBugXvIHB64fo4YcLv
OXI+0DE8iV0z42i6vEr22cihqBerC4RqV8Ra5mYsBUv/iNo+YeN0m38/wvOQLcoWNPNr3mmVNTmU
yV/faHbb+E/sGTpiG0p4VVbJ4hm8EnHIt4ZAfD6TzLNDvKH5iAQIFEnwar/77BDNNQOH2W2hiuqi
lUnK/w5NZQBFc11Uf25fgc3uOstmEH/vXB3CY4LmYjdDumau1Y/J/dHjWtJk2pdYez/uokt8Mr6l
NqPjyZYLHu07up+7LVyt5I2rLTUL/eyLf+oc8kFedQhZnGU3rXQ520Ru3rQa9Ll3FvcLosx3d3gD
tr6MOD/o9DRXBHTvgbPpBMB/TpQ4eLg05SlDO80ZMT6OxiyPSWLXsWishacpKZ2Wbp99VuSLzzok
+L7fMokzdiSGkkA3magRFQjaCGlTFq72qcItspLRiy6LhcHKEheMiB3OZ2OvMG1dYGqslfz6O0hM
ZKyRzPLgxmEBpwEF6zDC3mWlo3kS0liUy0wS4XprAcn+C1ZIDX9s4tAjyLe04OOpu5f3P0t2kwQt
2DKVpSBW0fXjNQ+7YOdhTQAdUk3wlYOFP/upyTTOEL2l+/OsE7bVFWqZWQPH4QDv05KRVGEUUlFe
4LbWiCcSrlRJv/s3pLVPMx5QRo1DqeF+Vkqa7rLZhl4SQ7FAsPp/7YYUdYQCps6xayPmWHwBbftg
qwq+ZxnY7MuTq20oqkowhTaxC6Adu4uCujgP6ntjtWVV6PLJbfCpKA4Cy+mArILSBw3zb25AmD3q
E0ngvfQI3we7ZZ/5pxVASMi+cFdzTkydELXJ/sFT7uLlTmLIMF859eTsU7nKAQuXmhYNAihJJ4Q4
hZB6rDX7I/6Lv0zjl0Vpto2zyxI0U6/udqkMfoLMfKElbHd4tgCN5/rlkrIoYqhIGMNIH7UQdZ70
5vZDZCgfzxyPmW5xcuiUk7uYJKXK9709q47JfMLItE9QRfpumaWboM+/Pfq66K4cVlcxRgruVdHJ
qzdfSIi6FItWkiYNw2ZrDmkRAzybKZ2TNd9e1xRO6jBWMclegJC6AYnN4z0fbWPB2WoZS1rFP8lA
vm9kF7grJv3QFG93Q+BsRToi78/x2UW5tCPhy150JW1inMFbCGBB9qyzrwvzsUzoWYcdbc73qPIf
Isfylb6+8Pv4SxlGiRWzs576NngXsLI8BDEdaeYga/+sCpRGpeEOtRlSsb/khi01Ye/umyS7n4/0
rJkTwlAbL0c3NwbYP7UGlseKK6DzRzbyoqaLXdeBk8WEfyUTiBzRKiVEWB0J16QHOQxabQ+oUrVh
rdNLG0auZSZL15U0uVYrpDNsn2+b8RatHdTXB3uHg4LMu0SCZFwVK1+EDf/KklnZNDbCk7CHGR7Z
Xbwa6rpx8UI03W/ZJq6ei2XbwumU3Uoi2EirXmYBF3qhSzfpJFFerckemI3W6i5XCodHaKCkxVqK
eRa0D9J/MbR2bKOXnnzeHE9dAVSsuXXYXNaxLnqfg9UrcZ+a5aD6/eEbEKUIPeSb0RhR2oxFUAYl
jd4W7rbUdV41g4FXC9Z3mMzyaL8YJWz5dfFgjpj+rbAXbjCwgqEeJnQXVHcKZ42ll0Q1HwOIN3fi
y+2qADZvJ/rpoX5udJldoREk++0pUVb6bqHht0QjWz4Um8SDc9dANWDoYl6iDShlAWN4U1FQFQSI
NhTfkIaApR1GZluCW3Ou0jGKAHAzCavCiCuiCA3+xIzOSMwqswe5Qq0xrwZN3TrRv7Lhz0pbDhEc
I0a5hU5SfSHCbSTlSTQhYnI+HS7NsAZ92GzhE/K3hWms4kWHk7a+klCsjmHgWAQB/eooZ2IL7h3J
tvbQ5BAYZ4gh8jK0VpIEqa2SE6JcugGi2RZOaFp2zrTh0hEfoHUXt/DrcwKvUPWRJjPZ37/grYo0
ETveHBMl6FP9xz9Le1dtMDZBD6+o0ul3TiYZyOegFuLpIhj3WiNIwP90GgSvO5Im0hbgOmMS45/b
PxWXTPoDqO+mizrvOq3kBDV80vmEaL2Hu//9RuO0t5XVc4YfahzAB7xwNDgp7SJdmof2FAahvDGy
ZuNpB7PGtbIQMDVWJHK5ihvUqPAC2VJ5iOr5ZBSBEs0cQL/4GTGWTVPRBSldjulJ2zhxjZJ8pBbT
PQPBavk9M5QR8FVYUyF9R/uJiKhRfDmOmCO1W8F7BoLpTQ1LCm1bCypHuSP/x9/i62bMjqglcIIR
D3cxky/c2uTfPopYdM0EDzKekhAXePf3LHbwUxuBPQxvbn8A+9CRoz4IyqaVzy0eiBCRARtEy/VA
rUB1kvrEbY+AuwAfPKEEww7mOjHcZNl+oWei5UuBtYx9FRdp0f1MHQWIXSpkF0tih/EIiW7bEz2H
cp3KPfAP+wiJquGtQF68B12GV1Q29fQEJ4s6OBlrP/PtKpaTIK5YO/EDNeGrW0ykk9Z3XsnaRTOG
h2y+B703Vd0+QeiMUH+sVN19cYlLMyy5NdDOPeBDmeml9rxwa/AhvViSOWnEbvGmfXJVGLxqTzUi
GBvZFRIvQv2QKkpGmYXc+kuO5wBLLv7HyezZkPZqp7iod7KAWVa+xaZ+mTMyqReZQ9O64cQJynAM
lz6uoKCh65UOWEzF9utg2bEFpfMTo1mocOGsgggfKAXPtjQuHoPQzvXHobvNmZiIKTdD5Ju0S9TT
Oxf3Hh+D0BTQbK8VcvMyp4sjdWHfkXon12mlNl3qorHpw/mm662N3Jzv2v7xyzRQiGwoavjCkSV0
cBuQNwKSSzx4Ftit0oIBgHmGFy80fi5y1I2exOQaNOvGly52h+2q606RJ1IzoPArM0A3JSMVrkFY
tXNPDZ0pRaEcqYBD8gqIV2v7TMOaxqJwxj4Wwp6zQc8U8UbIvBPgEAcfnJPJE5y1UV0Zw1RYWZr3
0g8q2EpQ1X8BUAmhUn7Z6IPKKVebkMpFMttUMp0v2BMjZljnNrZJkr+s/WvOJm3WWDAq+1uxW2rz
BfR+4RijQ8qv4oM/qG6ZDjpFGjUE/A7nn6JrLROR2pmbUUC/76k7+9nW/g0RaDc4yaba574z7O45
XEeDnB+Pn/v881TfuQ880TeXKGcu3UuY6wayJMvu/MnClrH+Jrhm434u+O5/zIizjgRrhDFhib29
jn4NoYkFm/qWICQgHo+83BmtiH0cb/RoXeKWUd9LekLKJtUPUTxkDe03WpTYGUqFywSnuG0UYMU2
VsbZPwffD4b+agJgXVa6rhG/l4oaZfCTcsWApLapyxYa01BvGtCSSVqBg56mComcT1p0NHGhS5xN
W/vgdDGBfLYFMqwO+fNSMqtSy+RpOZMV0u+OxvviaXDC7SQfgnHTqcjQfbX+9jCrbv+auI0SpOcV
e/RFq31slZCsJlarjsrLj6uSRR1MI9SypCWss1BDGG+kEk3iJZu3GE6u4qxKgplVSlftjEh72zqU
DBuDF14BArSWp5MR2STm4MsL2ruoBHY3v7nBH/dj0f44rkBlkOVUNLosEwVPuAf9wsQmF+uYJ4ft
noRnjwllUn30th1OcqEzeX5eRzgxzVKeFtBQjHTAL6KoXZrcyybWQYdiDBtYYM/EAFc4myyB5CsK
ICOil2uEAVU07WhpuUhY+y/vLhi3OqEYpKKroZjjv2aFr+1v9RqtHWLs9drWHWMK5ryKiE7PHiAu
b0cGasXAnONPHaI/iwp3GG4ACTZfFZiE3b9pOmICmmpPxD+tDhfGp4von7X8eRDSSUxDmmHGFE+y
VMKSwtXAi4TDy/2gRjado1kbHFzO5kOwO29/FAb1n7cmZTHZpQ7ZQID5qUYWNn7fy+lH6rG6szeE
qQxMQf2tywTuR4WerH+Iz3H1MWISqd/EtHRNnqGGq4qOVLdz2EV3o5eQ62QT4xTLgE15w6yf/+HL
jBZngtGYdZOgWSMyt+9FLS6y3r5tMx8K8XsxmFTidQTbS4+YemGctaJvZh7p5G6S0ADQphimJ/Z3
iRlr/9rX449iGmByPyMaSs/bTBwgeq9W2cyXk4sdTimwgGLFs97nx2zAqzR5YjnndP6AZs8CBSs+
6dmSgDBetvC8kVqpMK/tE0ieCbpLdnVt0Oh/2W2KDIG+HwCnhGg/Nl/G7mLNNMpnpX2BhhI8scum
XSEo/8TMWbJuhqktxHYwQ+W31cW43Cc4otSLBTLIEBGpXYJJtBhnZgGzfXPFkmtkNwbOEhKrFW36
d0yyn9j1kh0P74aNpg0RrtQI09kECI1mnmKSxMOLh46bo1Hp9UPG0bRlV1qZzIPVSf9qeyyi3Mpb
rzp4kb15IF+b2fS16vY63LIS3AahBjAKvyN9uLlJIyxk6R/fziuzYc6cf2K7czDqZ0Q2Ii/3d643
oIz+cGta8ewi/T1RX6eI4K8Aj8AatueJbsmXjZZdLtoHV8svrZ+m8jQ6d52BvDTGgHc/qlQInrD/
Hw1GJUUvaqfKVk3SOSeiBgCDlvmNH6hB9JwXyiidpdjy6xSpF4U8YRrPAjgbMOsEp0exZVNYbJ5g
w9jV5g+iOkOyVkr63WSareAExGf08wxWq+HdzMeSBaXYOZdO8T5+dG5/mtBReziE1rkdEOmdw6dQ
ftYFCKzkgx9emNapVcK00oXe/J+PfrOFktuz/7r/7qgKkVLEw6MnXBuXxRMExj5cDIVSM5wfXKZ0
YAXcf3rcFYOyL8v6cWG5P4uwYayC9fBpYq7PqTKwN7BQISqKkK03yIqGCe+nRt+UAoTHa7LBIUK3
Tlz1Bzg614y5bW0nyatgpIg7mmv3kKNagHx36SjzD8wp+wU7raxSJvSV+9Jo71ON0+qdrhnMYbDQ
t3Ztgxwap+e2HludN6OV5wu3YLjXSe+L0l2raXOkn0vo+edimKXm5EnPtfXv8DgdBPcbKSCTKsH+
OPtB5O2bscilEG/+S6o5fWz6sPf0C7EwT8hPkotiEAEP4Nhe9pzUyXsBnR9uhamKcvwU4IfDdaiu
3lVFmbOoHFoLaYvjG32Tce41lQmjW3mh5H1jRzaeBW7Xh+2+qsDyPBJEbKl4ZIHw6eV6q5s4VsbZ
LxveLwTDz0c4NeytqBmeXn4atmtlAGIIiuab4QermtKs/JN4wTUD4rvRTT4e09JP3ibqjUWeFVDS
4dhp3owRxCI9i9gAVfJSwsMIdSgk5ORZiEHoqpTbPJzlNpJ39AFkd0glIuy9/pIDv2zWRIhD/D69
A2EPJQsStRnP1bTNmr2KEJx36IZuJtKMKIEfxMYgdJRz+O1wCunkgbtwAWbw2878c3xS19LUYkvF
QENb/0xRSjmGOiMgShPjWus4LGpE0H1lq5KCErPq7Cqp6E9kVqmwbXbzguorUEQtPqSKMxixLOIc
HdvrswhvAAbko4C87v2ar45s/Z9tp76Km+/DxVa2YatUnIFkof74bW/IU02AIXGQsthJUq9i2tiy
+W9Hbe4FmsgM78NhQgtVlksO3DZJ/BjdZ5/+kV1vUJEIKtQe+GOCMujuXmILYk/PBY48GYFESXks
S51yn7JHQXaorWE3YN4wgtfCauqkNdHlZlfxXufM15S8XZj/VfxTbminc7accA0oVqbn9pWYvaks
OVw2GvxI0WeFOgxzPQdQcIoqvohzkzrtfCfsvK/F0Uocx0E203wXN86z1S/+2eZ8cCoZbZptffaz
DV06K1/vGlW77x7SZpdg378lFeSTb3UQz8rQwtsBdPoVcoIAEFnUy7ZdtP9datTFCffpkPaQh3iJ
89yfaEYMUoSzYR+iqZj6o6pYzMDqEWfjc0jDL+XVNvBQy54HjyaY8NY9D1mTKdBIWgb/8cMxZ5zh
xnmHABECM8LrQp3lx5sx3Ql3MooCZyAKtpmRpWxZFO/HfIq/JLzUhQwqRKuEPlaa8tKI4P5veWsO
2tuCcPE1HWxghRir8e0UZxdAYKz/FJA52aQKD30/21fHDAhjDDfiKW/zdeAO9isXLmfgoM7bNWap
zsOGjzm9DWU/IZiN83a5Ou/AqTsRsQqVkM1We5nVew+P3bzOGXXCjLTV9MzUffdJzKK3BunmCqiN
Ow+VC11mjT1sJ+Uv1TKjMD2Drb3dcNiYnF26XFZTnD8ukmRu+csCA9fdpGFxAIOvarShmuMrJU6C
jTNsX9hLq1gYxyt6xZjdp6S66vovCDetakctMbaGgiESkZUfT5x9Oh/fQBV4lTtMqQNQZO4DE98A
0LxH+lk5zQ+axyklrU9osAnvrjN0eNB6ln4PUIxisUZhERmMkZcPzgml0Kcu6EMfv3LG2wLbJarz
PTaZHqkaWR7pk7K0mEHSP8HwUxmekcX3D9eXSvlKOtMEB8bITgGdThPamMQ+GKVvU/8cazcL9B/1
hEp4g0/PPf9xfYZPcYe4/iewt56Wsbe4QTZWYzsbNRnQX8OZN9e4nZWRKeITjrZUPHNAOPbjROwk
FQong9q1NeNS0J5hLLA+KnSfr8LUmFMZa49XHIxHm9PnC2v8jQPEiC444k9WVKTBqJa109RMaKC7
vc2MY3j4uRyf5sonYbPyJbqBmxBbpKcvCRS2Y3sVrCNi6tU09LMphQ7QgBzpPitcYDzYoatTNvj2
94tPSHueTGc8OmMw0q+Tns44C/yyZWWYehxmg8GqefyejPg5rvlqFH0RJBiZPU+psPvidHyPRqqX
ODCBeOQkaEd+gLLQq6kYUcHbVSCWcmRQ2h3F2qJ4CYLmIoBpqaqoKS7FwV6B2UiRMGqPbEonmCHc
Rhe8GrSqUWc1eFlIOvfTHC26Bs1CIgoNDL4DT4UGUwVqjSrIA8rdhMoE+AN/a8L3HKQA51UigBHl
m3ri/eFj5cKIM/WMkBovNJpHbxGR5MiKz1bIvo0Gb1dcMMZKWhWGpuPdXOO63pVBDSqSwJom6pSX
d11wy+BbgsI7yqoeqBjYg2muPzRMyVLmPgXDFjgAnd63w8JSMyJvrSiiYvBseC8PYE7p3DpSEva9
fq8STuE+/pPNLw9BqXJrFffLZNFtQ2BXD8qptLISnNeDnQPdKjubhTEW92GrbltE4Ef1tJRGxk8K
8CnTj5iDhro1SN0sFuN1NUYVxA5090JworQ/SPH9hcGs6IER8BoC5cP0FuPqRUbCrPl9+jnSW32h
6ehg58mc+cdfkD+gec2sgcYHNJedghqAfHlQbO6MuL/bRD5ztLYSOnChrRa4WJS/pRBxJSamVm2W
RwJqwZtgCKljo6LJB4+X+CUPJHyEU7Wu4Ea7nxX47BCjDcCaTyfUaS6ZkODdJDDBpDO4GSb02yW5
l6roHkacFTP5+GOlw2i4+fVGVeUjHlRHTftXNU7blLxT8GFUNZfvjPhhOs6wbKe2MG/82JZP1WyV
lA2CkuyQXOA/vEJeb5Z532wspqut/gX8oH5u0zmZGscZ5oOjTZ8rrVcmliCE0sD9lZNUcU4+A6lD
wvUcI7IHZeC0U4HKByYzx3aZtAjn/hrtBPTrpYHABBKjzVk+KClVXHjbyZcyC/sq55FzShxoMe0c
xvtJ5XMxOtxT9Xw6zUp7cUtxYfnRbRLzHvFH+XjV1geazrZgpyLaN4lbRBgGHrYOzi7l05d5b3Su
9bLEYPS7ZwNswAh65pNFO0T3yG2rtv28PYzGJDz+QCJEyTPMmKRG7gVETjSc+t1Uh2kPaoQx1EfC
1s5tjUASaps5IKp4UFvVlCGZxyTBYWpaX79tCSR4HC0gEoS7Ms4EGw8gfxtYvdyYRgBtMwjb9TF2
o5bRFJNL3G2HTxBQDiHGvd6zvrZUcLNXt/dSbtjRpKhkIIcd9nL4KGx1VSHIoXjorsAvUDQQo/F0
p5IXJLbnIQ36+ovn+34+as4MyZjOoZ10W2IerjCjiSdJBDTCkLj0//p7rSkUVqaHPlr7AYn7JUrj
oOTNLmZxfjHJu+NHcJTejYKYMyX0cVO6X2f3g/VqFx6nIKJFD6vvtURYeZWcOKj8D5izKfX7YqnF
7Uj4xJiNKev4PLPIscVsq/bmuLJqvirjHDRnCIQuYfd1PKp4rKhRDLPRUlUdraI6kkMWRB96Fk51
3gay1RdCF5lDkPdct7IcPuQ0q0D/0rbQ8E7wVVhRkJmsfnOuN95wHU6dRALbtzZxomsxESyrb3aY
/ONXZ4NTe2hyqprdSc6zF9QpCW+gmTyxmq//peS0YRLRAL1D3Fgh8B+kIXaszC3YdhRiQhatSRJh
zxR39fPUa88Q1kQbn1Bf1LyIiiVs/6hnztmfATa1GdCqP5P/YUJQO2JjDtNggrUY7PbyEFp4PtpC
BgBM8jJ9agCkKnAJelUBpvG4V2UHYd8w4LuE+DgKTlnVPKENyHuiXESb77ticipv3vSJ0ND20Ccy
p1fyk0MRneG0UkjXIcKolLqX0cqgLHDSfAI5tqNBTWsvRyehyLGkAmje5kQSIIhqvyOaqVeaexJa
QZwU8omE5kwyCI6IlfGIh2l3r3w05ykYmj17Ns0/b2hKG8xnmwgzSwbap+9aOahpb5ZUzxVtmWdR
2eXsd76I0n7swGcLFrPuzyT843O7s7RQClLW8D82RuG3MN6kTsNdGAJdQN79OViPrykh+afwvfcm
fHD4OMbb0bLh0LGx/87m0bfdpoms+8FMOzQIqqb4uhqGuyg1gAdBr/fMqUGOOlNRT0zW6LIRXN4y
fcEUll+qYE8av4l/0Lne8x87WMSVlawK7sYdwClmDjPt6fXSRTuQeqODuqZle6tzJSPmPu2BAvgN
yi2PMDgb+JhfJsvCnJMoudBhw2SglYEHU9JebdbqC0cl4NBk5KRv5bk3UFKx2l5c9UCxSxQoDgbL
i+/gamWUDx8o8wN1+ZmRXwQadJx1B1TmIwjb/4eRDGRe92uRjFeB0MnUl+u0tslSPWkLAA87ojWL
MMPTlIxLP4Y2+BFyshiYC/wA/u9V9nq6HTPPrDaKweIe7BpXSVHCwIfqskSLqsWBp/dTQ8RdHihT
yg+TE4Hd/IxJI7hzAoNdcUrxcj7SGIS7punGdI/YsdFgAJQYttywXxztTlAMf607qOVyq+sU0FdX
ya5CpOCnc+8RcIG07jvzOYehREH42dEQUv7TKsFu0wlw8T3RiEOOctg0ehy5DoBPnV1JieupGzkf
fb+MoJdACp270UYVbz2Eq2p1mRWJ7nd9GwnufZbCoQKEssUXkOd5CpFpHxOKO+65LilYpOYLpfep
tkdGVB5itnl1GbbJOlmgbEfz5tbw4Gs0zmv1Tkgh7KRvPp1LfQ9v6Q3OxJd7z4/K433fHt83iFkB
Pe28Zpjvgibv4kVeZUC/WuWqCYGbZEhwCSdCCU8ZOpNVtG+iaSsqGuLGvsLr0tZYNLNRZHwh1g5q
JSLKtLnhuu0TH82jPTQ1/hMKN1Bd24wTFVkjNUFfG1yuQEg+reeZgNnZKE64u79HppGk6KaT3VbR
D/MTGmLRH4xYAnoP/tE7prC4H/m25xkCGiBS70HYbs0GBu4Rbpp7qv/79VRsJo31ByaismY48key
qgExim9Mm+KBa5SeRDb/45WJvG74+bLuOUBYSBJ7HCRFp0424jzUZQn6N+UvhUyaZaqPj49nngxa
Wxz63LWg2jGL1AopZn+q+H6WF3kxHnngoZHDoGA9bHOITiAJLhvYh2l0xb3b7Cqf2OLHeaAHoYp2
OcEbY7Uqq+WYsf0baTl4LUXDWHw8dyGcFH9uZnroZC3AnzPaQh+8/zvXA09g6aijnu4iA+7uuQyO
9LHvjxu+cgyHmRqbh3112DYMzrFDGO0WmFJA1LqqCxrU2A/8AP9L6dS4rdNIFIU4kSRm1SeXe5o5
n8QVYtx/DymdP3RQXzuT4q7StO7XCQSGk2wHuMy7jgYfoeloYOz8vxFiMpwkf/EvnkSR+jEQDqOi
2RUYDy6ovu9TMD49XoOo1uvQO4Kdyt0/xIhgvv6uAedmkbZTqZIGyXjnFE+0FPgkMXJsJZrq1Mmf
iheBjFc43dhc5b12ofgCuyvaJbSa5WFdkTRA4Gy1Jkf8Y2IEkH0jlhPWwt10mGTFrwbCRkyQ79xb
rEC4SlOkniTNZFHY+w/snXOm0uk3lz3DGnMphdJEOOuv/hoyWLAuZpms9aJKYaJoPv9gveqmsfj+
5g2pHux7O6lNwfwhvjF1xTUHdMsXQrXSPOTpjfAm/roqrc7BlccJRHUz5mMS5QDaUpL4JCfrtb+G
bNWYn+LlRD+ic5HJCRiM7+8Wehm3q0PYbnkr28dDZTKIzxCAzrEtENQaH+7Awf7dSUaOzVT+M+N4
srXG5/2JBOW+QjbShkjICZaknZFoccgvTHPm+Fk8TmOdm+9PbosRCFpiWbz2LTh5mRItYyYpgP/b
JIa4pKMN6wzXX0d0aVRCKUTD/fPp2Ys8WPrQMg4i58CkzC/uiCYZ+aNZgNM9k5bWeTlgtx/gXf3v
0Tqz+n1XRHKB/CkCrTPqhlSYvKJY7e3dPs7U1hbPi8OHeNWBEofAgDWu3fYby5FfhzwA/GeivHZf
WwsUUzN+T59OayqXH3ws69bJYuEP4O+VWgV13BJDrFw/wYumP1j1AnvkQCQB1JpIKCqfxGEXUNAk
n2+CAMVJ/iTZMDw2LRXNixtBMwlDlxH7g5OGw8PIZfNj2LhxcbHI3E6eMZVOpuQT2EaH1jTTjxOb
yowZIJULGkFgKt/qEEnk+C/U0EOOlGYkyHICEVIMc6OHZ5o8Zvc/fU0FUhGLxX+eqBKK5No3DL2N
2N7VX3LpD1FuM1tY7wON/QgtwkfS3Q0UMm9gysMut6vR2wtaXowWmSVhaVvzq/lhWbv9TEWmOKSX
rwRKuCMJ5zBT0CN7dswGBR8F3rrdmKmSQMrhyqiOXtroET+3DzEF/nXrnXcMOjneya5e9gPoJ24K
8BlItccnnMIsKbhUqNEb/JzKa6WGGUTrXNg3D0YoHdP+YDrQkWVPT05uY4kvTNO9Rc3S/LLlthz6
AHXQuo3iFAYwo3M3b+IqmQe0jTlslIYUiA478WW6doLHJqcphpoaDuJZR5DHBphN2P6g/ZL9GMgl
c2oLBusn0bpCvS4hKLBwKjYWVXPEovgHgmMOsZ5JXSK15Q9eKonRvGUI+W4CffpWM94FuFUFFflY
N4wSvF7qlLBdEuNNLPByBstrciodH2e6anqX2Mtv71EtlkBuZ37KavhHfwWZg28Si7v/m5gZMmVK
spKAZ1uxf9aqzh95KcFX/XMEe8cUXHuo7ACG+59fIfEFtL/ODRhI8PRHRaL5KSnzMoXwCyoS8ksv
vNB4IqVAq0qHAUwM1IF2aIncaC/t43uZOW6WoLTOzfhoLhHH7Az890GiC8fpdfaX+o+UgvZc2Bsf
MWAqlKxKIna9ysnEYEZdvDs71NBlEgioY0XZbDvDbCG26Lx1dlo0pmUb99Hygt9GGERIoILP4Wh4
8hsDJSdNLEodFota+CJ4oYpGxAZiKql5OCp5QaTxRWae94rE+XlRwacs1I6yk0GNA3sbphanfuGx
o5K8BWGHzqp8NbkVT1e0mi4sfzx1G66RBdBoqJe8bGaw2VeRbkAk7YhWCrl1mxhFSTSIfpntnMau
lgePrCQLZHtmWl/YdIwnohDeYxjFBtlRAANL3h1oCHVBRHLjgNpe5Nm5doHT2aYqJ7gZW8EIr632
RCWHHTbitVBqMnLeIhW2903poLH0a1g1lXQJXTQDdVUrmGnZeGWWcnRLVGZ7+4KENfvBMySuQNV2
Yd+3UlBlX/1G1rH/eptzgkPel8pjzXXfkk6OhWzQWk7rtjBkqf922fHWGCypfuckv0ynuLj5pzEp
Mb+TyqOr4LqVY/ekB0MwB58fyudqhM99NhZpC0oshclYpTZNDmsJEyYB0G465cP84DsayP90JkUe
OqAjwg1PhwPA6xey8ZsJkOnfoNOg2iVsr3sRnmE4E/Ven4c+8RvzEgCniGZlZR6QNqYcDR/14fmE
flQX1t7c7/tDdeAVt9lPLca7Su/4VympcGvjyefS7m0OHqT0YFyshFPdXB9qmrUWF7jvnFnM3C2Y
Y2/J1+4WIUpVzCc8IAZ7ajSwkYxCblwF2zyp0lfwxl799n/0DYtNkkkfqBuLeT7qYEcxdpma2TVt
mBEWgvkjbedlBWvaISk+C/c82rhwePO2/G0ZfDp6rq/k3poRNQ/8BQpdOj1j2z9Sob+SaLcKxpqC
HphL0Uqy8jOCydjESIn0WszA08VJLSJIs5UtlMDSgeYJXppudlSL95C5I0aFco4CLM5lZKqtJgOb
DX9oG/XlR0SPZoW2M6spoq4xIF1iqZLda9BxfeMusPqF4Ahbs9SdZ+DckIoqLahTQnIDkRMON2Gt
pD8GoirlN1tTUAJB/EBnxsDoUJHPdLpx4lPJCD54PptUzvtczDg4twaQRhWye1A5hH+zbRs628x5
9sqgJdQHcgKH7T/01C2mzItKfPjxx1lmkiCzyi/NPE3MNP3b7aRl5EoDAbxnrNRu0WZA59cXcOQm
x3ft9X8qPgn5P9aX0ZaNwV5t/L7ZNW7Ho+fz3AS2+198eJGbMht6KXEmgsylZjl+WwgYC+62BnGH
UPwdSiND4VVB2ZheWVWpKWfzoLU1vTGkImY4eYMcd2W28VvMXgzCoOQQNyZMC6iFUZRqKQW5kQPf
e5Cf6Le2RHp05KdeMWS97edZoJ4SqXbwr2Or00d/fcc4OI0K5E5lAzotMQWfCGVCEZBGaWq1K3mU
lzKOOPIhPqHD/RLOz81xdDQi3WDnpv5rIaGLWSx76/BTVyemAMDfWtxa9bBveu0B48TVI6nZyHq7
9uSia/sOAQ57eAM0NbNy1j7J8tCTmDJCuJP12Dujy9LlxzzF0/N58nU2dJi5Ak+Xn8JAGD/febVN
1+3FhMRDiJQ+1ksb+WOrk6uLexMkDwQwg/tRL6ZkXRwUQIZgJJR9yQXCo5OGzjIZGU+UY/rDGexJ
sbz2wiMVnG8iZD8lXqQ6nG/V81j05MMe4cgu/VLA/Z+uItHQmusL6g+WxSBdOdEGb1+fu9N6u4mA
64vn1sn4ByMHDuX4+MYnDIL1f+XOiqKTK8mgjBFwEIQbmLd8jjvjw8ipRUyXEMyGwoEu7N4ekc6/
cqbSqygeX8izGmG5n6LvXpkpP7xm1tAymGm+gbEY78XdkxD9L74u9aKCGf4E4P3cKzEib7rKeO+B
Y/O3He+SxTgVZHSplxjOWuzGtmFGznSGoXwshiEYTY6eaNU2tv/iJ4jgZ72EcUwzIBgEUOcX9teU
uLUFLlVX9mGU5xRljzkKwAS8WKFNdNr+vy9mo1YxnjCO0eWC3NTtWvhzQCFj9EyonIMSCq51FPBl
WJFxjyRj5hZowRf5R7HWt4XF9k8YigQNZgUwbksIjymI9xwaeQe6gU0+ZBjU7Ylh7WxfFsWIcTEE
O6+pNk3bAwzaBo88FzinTtbpb0duIEF+TwE7u3XWMK6U3urCxFvXXBpDXpVbqsfzbTbt9vJ6A8OA
aQ3l2HNxMWD30+xhp6Iq/cnU4WeAmrvpSw5DDZd9BoAlm7SGl1MAxr7GpXOFexbh2tjuhVCUfqwu
9ZTeWQzfdiDrS8tKhdO1BYPG+Hnfw8uawVNIlwHg2C0AYTFC6/E+LGYURg0hNXo0G/O0973HlLQ/
IbK/W4YzCXta62lUBwGFiuLWuVFbnzZ/SbPwEswzD+eyxUux3RtMTg8PvXKIAmHtMLZwk7UXAIIu
O0IjF4Up5U6Cx6ZsTagbE5RK4s2j2+OOB4dSRzub5fRvBWeILpMSzx1ZZchi4VtkTYwgnCOGU6KC
C0td7r5bTmw1pNOBaKp3hLjZqdJP8BmY3wjEhCSD6FSUjGKOHirC8lYhyBeS8Oo/rw8Z68fA3sul
8CQexU1L3QY+dgB4Uz+pDx61NGbFk5AwUc+/rZOLiF5v1y7AEVo6PMU6jDYi5jRZKO+ior4Y4y09
RJBuscPHb3I/NzIE/KlVMC9ER4eqdJ1XTUeBmWu17q6F6lji0coAlY/umGXHsUhcIpAI6bc3aDU6
4lluFYK90Z+xN87vqpl/3XtYUOyxTwWIWaY3ybK7K5nSvIER17uH+BZ7f/G5tF0Oy0yhINvDaN7X
Bq/Qo6vvlCL0t1848iZNp0ECC6bVZYeqiQrBoFo2AOd7W3mp5Colsw7OVZri/6Xn+xg39UmTbC4k
11wRtCObDMlhF391+43AZgpZkiYxlOFaDw+81Eg5EdUxAwx4VhYqifk8oAUgTSmbOBK+Y1BF1vSq
EINdK2BTOq3eLxJ0oteYDNFn/ZtPEXFBmpB6+UUKoU/cPPVT8PiR65fwIXubv5AABRqwi3NQZuEP
xM6JuGKfUnRD3+KUfMYbzvvYkapywxeA8qfuJKsb6iMXuDVSnNqqMQhOz4k6o4VeZ2gYBXtDSkN8
knIlI/gftuulY02v+pL/za6tzeChLOAzq+3kBAfmHqu3aMGup99SV56QyBGv9/KVbzxrpkQ1DhwK
7KigTjP90utpKAtm2UerauD9XR2u+YQhSc5/D31viPR4r3JYNATCc5zgAHiY+jxAwy4qz3MSQJR4
OV0POXM8eriyQn51lrtEnjJPLWPB5yFMSXr6WPavGjluEfhrGW2HCP2UhTNEWi3d7ke4UuTUkhIU
iqNMMqiq76uPiZgcTrhafbAsLLLVHLUBe44GOPhGWcJPlz11+C8ctMOZ1rW408CDL5SJHQvE9kJ0
uwUmn+e8LcE14wSG2gjkfe+AdA2Lj0bTrRhOJZuF0XsvPui5zKM/TaO3JGYxl4Vqzany8oPpSfiF
xiQpCTj7xi7p5Ro/j4/2kXNSREDQgGL/YB0xPWLExofqcUCyJDsuEnP72bWLTAuMMYXGpWy4+UGf
tYwA5dkXECbRZknW7Tkyiq/STgonEifkcRZlWnUJfinWeLD2P9wLAbz2WfR5Nd6AujId532gZnNs
bZ4dqyV6+Ju5iZoRnXtEvun55JknBNVhBAIbekwD6junsiI7qPxIc80ASg0fXRjt9V1Tdf7qZQqI
7KuKRn/KqIlH2/6MPQ3joRd6aHlWMYbzU2qvVcm2NU8y4/xQxAwO0PqjeecCV09txULVj4cFWM49
UbFzWkqNkhZZvz0QjdcFIHIlGRcmsLYA9wh2a4fK21TjCCArGxJvsxbQwTVQMpn9ihH1xRraYCGH
hB/16E8Vi5SYGOsRP8DDUVu6Uop9mO8z2CrDtO4pSjONHqUyTW9wnYY83YGHDw5f3YOHXZAWSMmN
9kC6Wc3U50qkyALNtqNG9uQrc4uNKa8cgpvvVEJej1eypbWPuJzHK0fmn9PDjBahYVbTh9rgO+Ny
hpHuQxa85c+zcMi1qY0D1fX50KhXo85dMPoLvToM+3oOLkltcTr+jRApqs1Augxx+kzho8Q2SiVz
ZCG8H8eOp2q48Z+UVaXG7naMBGovg/A58DlF5kfl6pAQsXwvMDBIF1cCc0N/vaIMsVrtUnFFfDdI
woBfMMrdH3QihknxvG36Vn35SI/sCjh6X0SRiU1mvL9Ra0rbn7Yc6KOdgf5uKwDeB7IOAR7Yc7Po
umKZYP6vwFOIzQdruvCFzvQEHouvlXc7ZZ8h46fHdKePQQzNgUEAvME/NPwKWhitQtXK1HSkJI5d
VAMUsvZAKNMJYhujy9/D1P0UkPlN1xVTgRP1iAk0ffP2Cmp8S/8Hexo63LUDUUGL7GkrXvYtV3vG
yaeoZ+lHYfFKJdO0QWa+cf+wj7+3LCa+S7cy6KPSQb/LgqEqvahcWWm7G6I3Ny4E6n2RKTp2yXYk
jkLtdUTrmpnrptK2ygNVllF3wJXtsHLfiAX9bB5KBdtHrb40bc6VVaeeDgHs4c/9ygXP7TDRPbS5
7QM8SI7PZK4L2LX+SYx4c1zPZY35RMeSCModBnTuu9S9Z97xw1E7kaizx6MnwkEnqhDy1aYm+rgi
MJcpKowWsgjc1uL7x1X+8ak4OlY1V6NGdSm4savgMH1oRDY3YlsDlLcrM+KyVVW9uwOckwXJlJ7Y
hwo+e6XSV/4Pzi5sFrSbvGX+ZAtHhg36bRSffROlIeDdWsIBstRZFGmEbs1TvoQsCd45kuc/aj35
WBbEbCsR885f+MFxFdb/cysba0D8kyL7zp/BOSJxzaz2+vUYTW5SbXqe5fFZJeLXyItYJchnHoeX
Gk2F3jr1nsDnJXwEWj63DbDc1LBZHJI0xYVqNVjCKHZRs+7DP2mSmY6mFxymCkCmI2Nqv6t5be4f
6GE8yEpZYMBCnOugSmaMdqG/dAyUKnTkLzjFsAojPnG1Ww/AkaHEC3FFN0ApYlqEsYZBlMZb31wp
RCBfum0FG6yIZDrgoJpisLyJhSQOxnBErN8ZR7PwEDNOn1uDjFWml1HJklHPsXY9pmy1Psk5xs/o
a8bUeVara8cW/64W9e0YUZPiFgmZEiDwjLc6tIadq7F5cI3/Z6Tmv+Z3XEj1blapey6eIoELcg3T
Ds2uz95X3HARNeJ4Mva9Wi8fDhNfnImJsekSxKnhQ+MMmqHSG8j6dGSEsXvh/fGVOlBwl589CNfj
F05vWVW0AwtfS7AQ0akKRKFZZuLYyKLwEdRsihqMzO7MdGLqL+5NBW4+mG9HnZCi90QHujFrjiUb
izjB3uPq4/JvZVCFNIsSVJ6QOo5LkpEt9MIJ9BB9qJMpp8aTj8iNSlawOox3d5Z4cyFkMeSeFAD0
bobtyUfRNwRi2UIXBvqG3IM8t0yn14RRWvZiB23/WdBISVgBflllGFV6aou/OiFX32+PJ47/h4bZ
bcCnZ6HI65sTIMRng09Ydh6dvj6WZ5QJUJ54+1jAmHCmNv3yccPP+l6d6jHilF+j/0eMxmbhuNBu
rDlWnxWVC5nXuISZdnJ5Aqa8ePVyWxA7rOk72ptR0JWAj8cK3rVmhU5a1PcriO6fIOBSZnUiLlGu
OJXlNT8s+AP2GSoPHgoM1U7apfFTz9FZmvryhhmj0VJBzRvcMUUK82+peD6U0LFYfUR9/KFl9wAL
RPvJkm3Dp/Q4xo5qanvBpn0g0SigTCwGUyNlEy+9ojuAQcdUACFH+g/g1Y6CWpaP2Ah3evs9+guj
bg2pAe/jV1Rwzo/oZORSr0dtp5eJjXR3ndFsnYxPj3+LTbM+dDXi5dYexsUl9GfBB6SR0BRrefdx
jJwEUGNag9Q6hv4N4DH3u1wBROtZ7WTZzPhqzJeBHAeimRswmcbZF2hDZfH7Ei9JdmWdOBWG5tzD
7CrSLXzNP+k1jcFz/6HEYpIYYyYghr+xvSHZROaAx8ibkCH0mJTX97bTZ1QRyVW/WUyRasj6mr3f
LgNyxsIValEpj1LnZwusr3b/PtT23f/I0+6SRReds+4IaMLQayOtO1yi8QuJ6msvL+W0TD/OFnVo
WOjxY3iRU1jxHG1IBnemqkt7jrCkjQeMWUCTl+mhdvZBpVv5sNsEMbY6NX3kLhVc+4Zar4eGJmWe
Uv52Kuo4cJAyq9FU9oCowmWXVcdMxRpysN5CjHRr9GObUkkihrLhtTdPX26UuHHJ0LnOSrk6kJoL
RAXUHHDL4sqvoeFRVLqv6PoqokcCZvb9v4nnuON34E8BJjrEmkySGS4Eo6Q0jp/nIIi+bONZ6gFV
f/ZuH99KW8RGsBEsHPRLFvlInUdUi8AnpC8e+pPnYo9267B4TOaXxkl/Pt75Z1zekDoMhesY92sn
/51eFGwasJSY9qoRm4Y7fGt7+by+dbVNB5G5q6jVcTT4OW9DeSdSJoJtohLQswG2gf4T1K0SW+uk
e9+JL6n3hH3yZUBTS3tJsZQ2NX6d6oEpiXKZpjcmedjxeXLlksesZ8e5hOK6ncifSH4260KP0yZ5
d1EOExrCytCt+Ejj4PmZp7isuFKrgtywToFDAILI5euvD/xSxr4jZdy2R9ch1D/ESHBZl+5hTfTH
O9Cb6Gu65/rhhEI897jsE+uJbwOyPgEecczaNEd0gc3ZveqGW2xtsH6rgTO1NSh0hXThbjGHW6/r
KLd7+0na2ZO/DjcEcFQnqH9lSuirP7um5/I8STUpI9iq0XHJcBRTq1bBsSpou1U4Wsm+FJ6HQ0qx
lEGknfO1XAZoGVGgF1xXeIYnbGG3BuNEJca9R5znf+2sBtpvDj6khzbex8OLnO0EHArSllHoxz3V
rLSBUTIPxxDvTVjHqS1AUOqKqStTcfRuDI6v8tlK1fs5Cpy+bFWcgR6OvYZlmWXV0AAjuw2vTK1e
cHA2zkoHAinLBYYlFqJBNorzAHUMy/pBfNH/ICHCuoSotGjD2WQ+MwMdlmaGwakCp29wNGzwQ+QN
ngpnzQm7BdM2eloh7Nv0t9yCCQvr9GMQgkVe0swSbUI4Vgk4OQR/lNr2QEyGOMuT87Rb/JWc8280
r8WjbAtfortJZPzYuHj/6cKQhwzIwGPqmx8Qp4rsOn0KDT6tGsPVLNLsQHLtm4uHMhkk96q0RA1i
8Z9EflJohunoUd2oEi5azxAN+99rM0pGB5mYGgh1lCU1hkKeWz8MBpwQhNt9FlgT5zjiDU9jpNER
jAXHMF+amMW9YOXB0jYjOyPjil+MJe9NPTwaigAiPBONdoG4SVMYMfkwFuzITFPY8s4O9NOpAGka
pQV/Tw2gpn7UUB5Ccx3dMteorzb3/HxINd4Gx/YrSHRa9jqFs0k8nyUC+IKjS2djPjTF/Nn/tBEe
dNI2pSYf2C2NWyRW794pMjaDyxDu5LbfqgUqhVH0sPC3io3QX6EiyI2TkB34Pf0MhFtkFQIbh06b
wBGyEgHkQtMj2xJyetrypYNEOXK9soERn1tNuSMoEDRbGupqeu/ToJLNeWNRgnOwHJxcZ4/b3QAx
FOQ50wkWoXEaUoElw64R4EfXs+Nso2ZjrBKjKoFm5MgfVcBY1FMwanjUhw64IvkBE227BPcgSRH4
1IzivXZ6O9A/RAHudFKAMbuiN8BHNIeezajYlyf4NW2BrY679vkzEEZaXh9BhmcvVG9AiMupGC2I
0rrirr7D68Ur+hNhtgyNX7nqR7Y9mIIZaJalcb2jv2pwvbt7ntKYhXXFdJBPXuAYHb0KTBR26ke6
VBajISCdvwAaCfSXmLCoIdJmF4Kvy8v/T2zgNBU7SlHlEuc4eMCmAYz4GPf/IyOzKLlALMxkBIXA
HsBEBQ7WOkwMC+6bk0NTwHhqj1yqoXd4lS7Yt9xdxGtEZ1KExWiGFqPqO7O14mxdoIm42XP1T3un
v2Vu/kKYquoljciAmgdoUScYwdeVo+JcGQ8SJWn3d+J4sCc1emFXJq0v6w5QAEpm/PfJ7fWKxCHZ
LAcuta9+WgcupN++HKP6fWeJGlW+iECL55K761aPRNgQ/NsTIw6ydoDR1tXVhNalx9VIHU9PPKZf
/VCtEioCDInevDMbzIRk7Zzko5dTjoEVY/86g9Bz8A3uFhk5/KZRkDXuzY6BjPzQohcVF0ldUkBf
Vr/28cLLLw+bl/jlzkQSpkAXAKLELG2/qJjBlyS5zn7sLs3/P3qZ21OQpcja5B8n+h/gMJZyJP63
DfZj3/hk7VcPXjWrTDUokilreuj1GwtQTE29EWsCm4prg5tH/mCwhLrQPe/ZmzrCDWTfBNouB0kP
uxh+w5UuRBBbtreGSb48pejdMOQqOWx6lnjNtL8MPxcqmakw4lpx8pLlbh0oBcKNr26qgD2vEZL3
tG7P4HSCpo/h5/+sFCtrtqXPm2KechzmYqylVno85pTB9PEU0/9CGxCdJb5qlPB7KvXp41OBCG92
IIK4vBcptLa3jmLA7APOama35KVl0yapEBB9dFYBMdHXECa8VhYE4omPBacr4/iwpI8N+6PXflv8
oHS7IYCyUFvQo1ga6PwweIiS1gmMofXBvUEgKd5MJSkRbuWOHNKCOujtyIfn7cTNju0laoP21Jy1
UJcLUBh++tsExBmXjAOqUMFfZ0lkuyVYet3j9WrRtvrFbzTweO0D3lobVxgZqX35MW7OaUYbnRyn
ceu784O6HWvDSZwjLHFrJFVxtQeuFrLc17gLPHEHhlJqAJiIj09M0nw85lNA3IS/lfrUbcX++hoY
PpeHQX6vIeUfadkUldbHyb8lJMhsJPEoNGptLzLG75Fo3u3Ni5ojDJZCAFRJkG4TotqZsw7zlTM+
/Tu3uR/hzJU9TfFTT7DOrsSLTHRjrXH5wjlm2W9mTGji+zewdkyebcL3gkZ6VyZgpFbsFRrbhWrr
zqcbaOj0F5w/VASZIpZ20xk8z0/l8tfQ/vfnvcbESnK06K5A11h+p2NH8qpid0orpnJSqDC13/lS
UohzOq8fFYepo6Kzb1TGhlEONAYfYZ9FBKNjzuDqAOp24BvD34oGbx0xiad6R4zYt6NR/bZNX8fq
Eow8DshF9MjxCTwwVOr40ILLeyaOWq0447jAg0yA8hRhp8OcdU8D38kxxrMqRTLSchZjQeMT0V2j
KE8FOrZwxVS2c0jXlBqhdozsfA20cgwktvRocrCR9GTk6xZ1wIOpJpEe8hI089p5IHepmXM8kKgu
BIbYXztXl0fCm23r2C7D/E3kytJZUR5YH+QCnUOEn0KHTlkH4gQoERgCBb+/xdSrJ/zpd5a0JYaP
VRP7+EDlTrUv6QsRFyc1IoeIdDGB2+cXaxjcQ7o0maHYAS25/2y0Eu9wLHH/oC8Q45iXDNr4TIdc
WqY+bnVHZEI4qowWKo77BKtxCTYyEfsBTHvKNuBGZkE50InUtOkvLIlO+iIerC6XkV2RdC18GNjj
6j8ZUfloEpb5X1vc0J8hUyByySG33iQ3MlOwASEqkG5Qu3Qpep4WhgrP95LdVhMCvo/AYw2RDC+u
vKGzGDjY8Sk1xKnZPKhasc7x3v05FElPcPssAj3eOHHiUmGpzWTwXhxzIfoRa+gJHH0YnAwNG4me
rXObrPQ11PGybeEhCE6oBviwZGmGh8wI5kNz7MDuezHfPDdTrzZ0hRgpdzIzeLGVmdeZqqWto49Z
v1HyhkTkFa9uw8uFLJOtKxtl8oLJ0AkWufEM0mmFKYUKWr2oetLDkeFnP9tvk/xZJUTFVtirgNEn
S4RqIfLNVTkkm0aKfnbqMLW7fFOCocftdFkcWbt4M/LG8dLObqFrudRqPLqHMjwtu6klwbAH8Q2y
AOunufRLEN3NgYR/mAIg5BkqadtDupyog8D3WqBuRxA1bIiQQi/qVF+nKz80KgTKcLYynSAEqXJf
tyyMVEXg7ZGooqBPFSu6j594xmKE5ey7BNZvrq9yOp88b1zt1I0wABFJZ5ESBxVXZnHcrT8NAJUS
LQkS3eyLRtdwpnyURVaRp5XBLwHkjVbS2VlcSLgYBDRxiZaPwwjV77AIWOiFY5VCAC4AKWBkB+pa
d67qCQefXoaKhsSt01x2GntNh/7oqkXSSUTHuLsNnKTVHhaEj8F5qpMH7VEE/AK88M1ZpOohWTmj
Ry90cdr5mjSLuH2yMqSnc2KpiFXBiJaODt3lc+L/pCD4kdegB2HgsP1uZGSivfgtCLeb91ubPtLK
e6Yic1ffnaxD35vi3ssdOvaRuIcL9AFPJnd1YdgQxOiwLaWcCYTxSGH8T6/wq1oFq6NUdWO4++Bb
XrXoa8jfTRHZurzkio/6yMGjSfClBVTDn33XYJSH6u1p3Y5Tn8RrP/OhBMfCzg8soo0x7mhVCo50
kRMoeq/bESm9AZzcJMvYBiQ4hR7QrC99GnexRuhpCGIbqwOVbQuiPk+bjz/yJf5+dQ+ZV+gZwdcp
tgWlqL8Jpfu/He7e4XCxs7VoOTuE7ff20FKTgzu6g1jTuXpHOD/ia8kefGcSfgzU029fUQUhFq7u
M6i1aGt/OdkDTuFHYqoYQm7KT1iCrqiVAKzrpWZd24nvD3ta0HIyfM8o3yMJLGdN2a5Cj7yZZ76+
5RnxVcjhRB9fA8NrhDOsc4KI9czU2EPf1mGzy+rqnSXkzjMIgtjtFnCVl+LXn6rGMU1FPkUmVYeW
V6cg2/2q9jM/BMat2K14JkdJXERMwlSy4s6lCzTO6Xs/C1S6QbIzQiM6bXf96do/2pTIfKM4yGG5
oNc0XCedRMZF8rhNjBeo9morN0PZo4zlZyhw3X62yZCDyKd43y53+5eRX9TcM9YZ/rVuBew8Rk1V
scBropR3emR38ThRma9zYNlel+9s7WF2zMS92Rgq95f0/BTFulsEnhQSAsJKinAwHtL0Ep/CoyiM
kZcNzt8jk2YUvxj/Wmfij3v9/848jjd0hqzdUvBNMcLhuYIQhs0DWweNmr+u7yp48Z9lXHxOhT2X
QOgqbuXURn1nz9Rwn88ULA1+Qc4xhqAsrCClmWgQ5eEGkFvkQvdNMxuvKLGOAKQM2RhKDX2ISmUe
AkTWn1wgfUTC/1p9EvTRdzz8jTujNmJvPVJVOJGpRFti0hfuggpeVdKi0xTR048jiwwe1Y7TdBQ0
sUQF/SrFltr2RfwWlozcujD0Lnzb5WfNKIM1EzPOakb1zYHAnhryYr4N3PGl35BTCzg6dlRdv8ek
3gbl2prXOK0SynSQkIbGsK2u7cHHtMmIJv4hsJTXnFp6ZCp2CKgq/wUD8s60xAYZAZWSBjeWqi2g
wTlreNoqncfxM15bzfNtoJIlDSxWKx+ttOTFjCGJLilOPFDgD7ggF18uMYenGSJ8A+d80DlsJv+Y
c1FNxT35nKuXxwYVpXsXb1YGwPQjnO+e/eJzafmtPyrPMqyxU9gc6YFIuf+ito46W2DZu+yXZAJa
s9Xz/ZMTYHVXAC4DptrWkRdo8063/r4YmtpdryTJhnKfFD/QdeT5BWPFv1MKWJ2+pxhrWTApUF1L
O0ou/RdPwIJ+3EJDQp7SrgUtO0QSJhwna6a8W/IvK2OMaPszQwO/zjOv8YMXNMhByYh4Vv2ZSKei
jEn4HywYrxUCOy5Jiy6WszjsIxD5pvdH1/4d9/Lz27lm0xA7uLi28b3QZFbDPPB2mRoYxFZyjB9D
1OHA3goD9VZhbUq4quXQoEoy4PoglwGtRmkn6IXMT28vvGuekbH2vkg/PBiNXnYJ9XCx3ge1dhIO
i1snPXaqbD1rVg2qZVtUqFUx2z3yjjDyhlMN3/Pfu75tDbvMsxH4QEzMB1o96w9qDfIYLSFjFW1M
f+s0RKbZb+zNTLYU6zBB69ksFifqVeQiOTlw0s+VB4k5M1jpTIBwOqms05fBTLXxLPpA9f+lUVId
Q9Fa17hgilaDjg4uA8U1Ve0POuB7VZUHUr86IDfwXQy0aQLBxnihCmBoHlvDWPH8wlJx0FQTISSU
KibzwmDzU+Hd0nuJhpH4cCpAG4k432unNJwUC2JM5Dm5YKQtvvpulsdAv3VcFdNwhsqxtTHEEB2F
gL9HmoSg1g2KY8FW69WOWUi4Z/qEFb8m9+GTZ8Ul69mj9RKxkx+/wDE5/GWrMCPPFbLvr+OLVSQm
qpgLtCpvpBvMwUYNJClt8VRXTCDXvxCXJJ0lzaULBHWbgeuIjZqhh0kny0XtBFVOEi6TUWT2yWPl
Lewl0Edjgk369A/pR026THnx+ZIKdygaXEL/2+/Bqb4bT1raSum1X9XYtMkCw5L8/jEc2coyxm+V
haUcXh6C4kTJUUWYBiUqFtiL9A9I5nuUiz5p+LBh047TcomOyLzHBVkfq60feqLXV16ZTgy8QFxV
Ts2fn34JsFCT2umf1NmKGeYnxN443fN4mChhfO2FrV+E5rbAO6wCNgysAB36mOKzVGFqD7+KeMDJ
WoHtHYryWJ+h1RnOXpAtuXmT5jCSXXkwSBJw7OYZvMp1F4ZninPWhf/wBFlqxa33o/gCeF2ph+z2
jD/I5xp56nSzqmOoqMcL3xfyEvu1hBDco4HkWcLhcHACzAoBZQFuIqnkTWbZp3iPrIq5SXLrzpH8
VvrztoOXgPbhCZ1BbVIsZaWQHIoCqhtxwq0jQ8V9kZ0XAbLX3WLZ/YHVf0xVcUlzKYj1dtCLFzxo
CCDPkEX21/XUNrUyDKCW1RufN420PBU5rQS3YXbHblNYP84xt+L28NlXR8Ur8dNYP+6i0hMAwqqu
tEl+j0Oyuw+fwpRiZ14u6h2VtgLAPyVNmxcHNryaBhCjMhFCFLmKUuYUlqVyCvW6Uzy9HG9tzCOJ
tU5uUZrCClpYBzjJHQ576U65qM7ZQQBpkmTR/2uotTcb/rZFM5FvMdGjxYVFRXwlWmQH01sQ9ZwV
AEYKzgcQjwj0Y+/5+Ae1ST6nhU/YU+R5mrqwmxX3PheNp4Hoiy5hwrkIl4GT75NSBwEqyrwm6jQx
dJTB8SLqBDwU+EmiPK6ztR6Y1Kok/uPXyVSaIUGGr7EvItg2jIkNfiQv5B1cQA08IIA9RflXuRx6
k6ci3+Q0nTHyVDS0pvk6y3qDWb9MPCmAhX4bzg9CyOWXMuDxD9Dr876oTNpza8mxx/vrH2fOjcJB
3YHA/E1/Z5jeW4Ar5fuP7tn1EyM5RPqmJ5vmj8UP4uZM7JdFBDYKhHYUkBzY5FSgPZk8hJYil1eT
D6og8gdL8QxMjwCHCZZROvEJ9LmO5mLIVrMdTs+qIvkU1sENPazA4MDbimbFEUr+QbGpHwJhysIf
7byYw4cJC38Czl4kYE68T2t9eZ9CWtRB3sf9scfws1vAw5NC8UtzFMj1vTPfjipegGcdjHBkb1jG
IacwvUAGHdlVba7JzAJJrxkeTUG5NTQGYni63s/E8UeNV3mrMa4RHIMBBHrA17ge2qFNdeUUc0ne
sGJEJ77eCzwVtS9pg6KdIYFijU7r/qtF/29FP3NjMhhIASp3QzaHjkUXGzrzrpc51l0so+ygCMiq
PisGbXC/X0IpNhcGtSVQJyaMCCJvI5GdCr4O6xMDUiso2ofmDjM5ptt8zVpnWEHPF0P8rhmH3bb2
n0Fw7/iJMl8IXC2fRcIn8M8Ft/UPqnV5Dppz2NlKkXwWDl3RiWehKsauCbm9XtWJ+7QSgUw1UeIj
S01H1htnn+qKG7BM0KPTnuH7MX8ez0ZMsMvfJGXq3OCo6K6ssIw+hRHWEaxdSBXyY5RdEfRqf+3a
OcpVvps/QvLYsJRPqwgAq0WS+dRR/qPxwa/h0HTymF9kn3a0K/5zpbqx41Txv4LsRgoN/T+QVGvx
A8915KrcZlAbLFr6DK9a9Ffk33zGsLaMAld2oNC66IomYZuHah4kpcTTYPpMAX/5zmasQhQjkD7E
NYDoLq/GTzMV13b8+F4ela2REM3X6vM3y3DCQNfViPj9/5HLI8vgyu3ut6bm1/USqIktaqq2hCEf
bPiLN6fG8hp06weVvzNR6N7ugJ7czdv37B0hUiZyq7B3+JqMz7ZZGCF6cr4/Ss+dHLISfWLWNH+l
hJZakXDTASFenAjaQadoXsXF6IGGA5DyXVqURGujrMdMTqp6X9Tj3KLiQC7q7RFbqaa+cIL5xTfN
IDy15d05k+DhphpObgGuIC0j8fvnpIyjRTQwQ2eSx/H35GmjNY9IMwHWvo2lu9CbJVmBbR8WIltA
9WSVLdvco2BBrDJkG04THrZ71ewWNskzQox+3VmqLRp7xvUt0dtEsQw/w1uPRKA2ClITdWMF1vpZ
AGQzEYdPHafZf3GhpdBeaXwO+wHz5JLMcztKJSiMi8IMZrMDrsuVit4/uv8pXXUTA0UkObVxMpjy
1NdAMAtGnIEaGiFywPSPlhDRXEoMXbbY5W1sVDmXqhcjGLosVFMzqZxO0l+vorkmrNSTDNSDnZC0
jbkBiwLrnJGsxdc8SDgBQPbj29izYpWwyy3lC7a8kijp3o+yi9OtwElNoHNg3M+ZeKawxGZv7quB
CHjqAu/iubG6ktL/SJxL10jHAmWH3h9t7PxBp1qVWu7LxIzNKjFZZMoL8kHcEle2zl4UMMpMY9vx
eMNXa0bHzJII4mJo56BTFyyH0oygQzpdMNuX7V8rD4ivKEs/Qmcbbp4IIZlKgvp7DWuWT4WhXxsW
S7HD2k1k9AZnO/jR9bKV85mkvvxW2ITqiu1p3eu7E9GiXs1vk8ikutJDWWfoPZz0n4+dL6S7J/jk
yKY3QXnBMNs6KRPqEPHkOVz2Gf9437aw0C6x8ZVuUjJMc7lZg09Vfy+rdfbVeoRrKAqRA4mNMTtb
U7601j6LWWVpg62xyJzpK9sNVe4XDjgBNz6tdQTnuHpIroKnXIeFi1Q5KOIHYmADlZskd9lsciFD
iCwZn1JIcJs1a2pYs4xHOdS4LRRGd9GiegPYGapUInHPELN9QNRnWawCmVk7RbGKgdopdP6+xr1V
qc5a8rDk6+63bCFT5tOXbh7pzOCkn/00joKCOgkPGI7Vftda+ArFWdNOo0vpi60kbHyzu8qt891S
4N5InUQtVxXl1NObusYsy8J95bmKlDKO5Sj59DvVv6EFJliC5+/kygDKxpav7DfK7LjAOdzK65jW
qctC6AqUyVwoknPrKjff3a7/LYPvhDocRRLQ5vz9dxBTvQkME6Rgbv70TjR4cEEufnt5svbZc5dx
dI1hEPEOuIpXK/74fvBZIyYeXYowPNgWufiwVoqHzfzd+jmfNgl6IN2fhEIPM9V5HmSwVXgTjF7J
Z+yHLMPl3wnN7p9EyjmEsPHAA56xJDhw3SxpWUOaQ10/fERc7a9D6UP1etMyFfg5LREnwjY2orFu
jt3gka0E9l4fdPSfEEJ0v/Gq7wbLBc/LyOv/o0tAnDPZMsvRZE7Cnyp/6akhb0rMCK1OLkYwTRQQ
LC5vkt5bbUVkZ2u12MnWeOG7m5bYheA0pCm+MfR4wKcYv66MLEIt8jtnb83ELALyXpF2BIhWvfDf
rnrRfvxcypOqLpZq1IKLLOl3z868zJTLR3FfzikpyDiTt1MiuFGirfMZQob76DUjOmN8GPOammPD
LCvRxst1Z9AdM/uX7dMhpqHCWKF+nepLaLCuP6p0h7vpciQrjAZFjw+Cp3SwOxlY3UViLONVbX7l
aWPjwNRsdEQYUPX8v28asnH+MghihvJHYMdYuUTI3rCgXM745cB7yAz8mjoBQphq3+Jug+l3xyum
CSp7JHB60iYJbn9V+/yWc28qFvBkKC4gxy3TTGsPU+ucO59uC7M78l05IdT5zi0VM8HxpTtsmY5r
tPqulR53vfjDNcZgGJmOcmTBMAk2aAuuyrKKaq5DmEd9pmbKv9aMNiET2SItXCKT/Um9sTaKnCC0
tKBKqjSRwcrTnGTNujHREk7Z0SR2XvcvyJV6GtlNHzfGlUbdDFuZI3kAOGly4eHpa5UWEgrLMjo9
nMy0pP0jDMzCN9Yst+qZF9T+RCp1YeUaA4tgx1g7ltxRW3ISWqTQ9T4helLtT5O/bKj5RFFZp0So
2vwOD9KHj6RNfMgnOmU57DqrSvYzEsT+a1l4LflkUA0sNXMubbvp5PJxXVxjx29ynRCXlyvGEo+G
wCUB+72Td3VsFNiZ977BBM9KkbLfdcf2st2TbD5YJpLII/QX97mf7TyhWdN1innkujBVyyjyEgF+
qdRpd75v9+D1VeYOgeB9G7RvrfA149FjpVFg/8SZWq9CL3yajXijvJp6O/vqgM6vZjJc7f8XDRZS
dbQYkqjIa2Pfmku1vK2sda5VfAAPkrNAinXAW7rK5pj1tGHXiTraNBfzeD4LwbCerGapJVixou3n
1/xMImdNA9aK5SqOKokt2FmSz20Ov4Liy1eLilTWizVZMXMPEvNT2KI9zhi2rzvazCoB71BUUVhQ
Q6psjWZzPd1wVh+7sm+QRCf/ri4/rG6mSBwy5tEdp8rlCrukCKYfQ2CJkCVufqtdIJGZVH9mfxbB
9fwe5LTM1UgYcZGBJ1S/kKR8ITiGNYXvaLcs87GiQYcUHrpOBPzhUxHLoTaSUGLFhDhgPABG6Ge6
5hgqqIf7RuMcYAj+1I3R2PYoAIASXdd/OZd2uCsq4rNvihODEn74P0RWR4RljGOjNXNXI7UpV0rf
hD4wRzVZr4AeHQG56Eqey6LYXXI3PnKxtRs182gOdyh/XYCM01fVSseR/IN/sduWpoYDhHZtrnAB
u1LAoYpKa+RjTaTqmY5yqagTkq9q6wTFvOyTPkgMEz9ovSyKZDZgPeQ3caPujm8yspX7BOaQAkGW
o54Zm3lv+O3ti7ckHUeNbZB0lE1YwRKEv0bzVkuxERe8ZK3qhWKnlrtMsggi07E9l3jQmVhmuaeu
XZwJ49nlxg4fjSJWe5nZSrVxOBp0jYBVef608QjuHTQ0GuJg6/mBuLC5SKmMXS85fJSh48CT29ur
VnwjOoRrgMKuNxfDXvD8GoG0pv7QCzXZen2CZBh5+DzK90Q/om/YOxkDIFkOMKYlIQLyVS03Y/Ir
wTgvPbD7xqjvOAaufK1bWvbGbmrGOkFMb6QnBC8AW84kpCIZCBLRu3pReFUc4pWaA20wPnbUno/+
jL1poW/qfHt7KU76r+VrC+XD9brce8GSMHv2/ozpNWMFiWgilup2SQxoX+o8j082KxcmPZQYPR4M
nZtpV/vA2YcYtbvRVcTTJt0v2rH8y7JtZh4WOHC4W8a0pSx+2+TdbBbZxpX2AIqVNuZWA7yOkiqp
ew58PvbkkAfVGNMGa6D/GiEbwDw20Dgl4YOF+gx7B3LBsL0nOCw85ivf9ysmF+DATuMEIIuHktX4
V6N+ldSgnTpZViMfjDvHIVj9pZANQD/n8Buu4STuwtGAfXGl0CL1UdrKcU3TKI2elSTBP6WO708V
0GQRFnZq/LlOTUwJDM9ZXo4heidCWXTgo545mRfnoes0TAWqFMUpUOz93rvkYmEO/oa9vqA1ZpsN
1eDxX0oZe+OFZwTrAAgRMvZ86CSfYT1b55f77yhz+gYxNLTAo4n5945YDrZGAV1lC96v4lg099dj
JOgEMhLkEo1P2XjGVrmHQYgC9Fw8kNl1nKu00b0eAt9DTZ2uR4aCYNzPA86GtJCeua5jD9k+gcoC
A4qepRmpcjRRj6isI9M4wuY9ZMqr7S3U0sp5QCqdOfIZkZcZVRjfndIbnMb4ONWAjyvDR8DTRCv+
3cuNf4gu35N5LROtH8mCfGLoKcGbsHEJWadXOi5ao96cS2zsiv+ERBsi5m4AXShd/bDBqhgvVQMw
dT37mkbcugwW72AKuxs6vTyA/XnKAOBOa0WpAmeSETVI0mwy18wQS9vsT2BzExHiOD2XWwbXIlyr
lIECN099NfYXg9nSMyXQTz41LpcJ0bByJV9VNW/p+hD0puU7Q9n8xGz1BlJ4RvX/u5qzTDOvpOpu
eEzfhVzLL/TxyeUnBSCA3f/v9JS7E5CAyQ0NKUYtaX+KOXWA8DieQtgOv/W1bogIrGBSdcpqBOHe
P1gJY47naaDzyEpGGzTooFA2hnaVH6IY5WMdr5y9i5QNhDWpXkgEcoORGz3xFeeY66gykMvGRWlo
ermmiXIEXV6hy5IKzmF2Cs1FgO84NsvhBVE4z7dIGtSnB2FMglzF+0a0UJBww+4t4u2nMVwMkZHb
vz5hXLukLrbZaYee6Te+bF/jc6ryWX6VyQ9QnH75MMUGQUpNlD4AA+0D38Uj3U2fiJxcx/+svuHZ
uzB/JvNjS9LWBpybFHKfjqAPiOUkvphxMrYn3Shq5XFM4X5oXgweCXKQIrnqbTSVq/vmoNAPBiqz
EPrGNfxOhB9Xy2IRuBc4UztfRHuMZEZ094l+J7PCbhi/lF8U7Bjlh4DyHAmmda2NglTriW1rBLzG
rxHmU/jfQTq0eLcHWcnrbMztu4sGORA2lGt8gvFwlBuOPoqM6X/icuJfNCOODD+C2spi5IzDZ8jZ
N04mw8R0aNzyhRJtlPgxI0hb+EW/aS8Gmic0mR+d3zdQc5ynRPrS+Ic7+DAblajSjTGY99q6ioYU
IIHAYJeQulQRz+cGgG5p5YM7S7Eh+VCE5tDRBPghREb+a5+doRENZWuxLmyBmRk8diTEI9m377aO
26SfA0vFv3/X23dVN01EHCuzRn46kgQSOvrz70ZYZW1KlwLqy0gB2iMIJskvdfcvqF3eUHzAMhd6
Bobul+QJZMIJC0NXndwjjzZWhvypl79z8mF1YD4i/zdrSZoVWwln9zPRcbZLPz5WwIJW0booR9IL
eqMtkKZ2q5Ms+TMqc2jb5kAR9z9qIH6F/vOvqULDEGTcezalsopZdAS9C8+CtvL26ftMvDD+bwD9
FmPP8TZC3EvYnoul5cWS+6WItstZ8akSaEdsZUtmWefmdWwCI/oDKOY3WD8J+xTkUXi7U+FXyp5F
lccaC+i/SMviKM1fkEtO+HEymMSZqybuTbg33K3YnJw+cpP6ZC719AfEznsS+OUBsqbxMPbEV5dQ
QuD+0Sx60a6BmykXaODFGcwmb1DrjuYNbWmmd213E3XFUWJbFCp89zNyA/ICN2APfYhiw4PfKg2Y
Ik54YImLgjlB8YEY3edMg6E7xOxceRvwBXAFvZurqy30GVLg4n0wSrxe6hina9gsPw+QlkRjK4r/
viA7QWW7GPgRKQ0scVTdddTh2NkjBA90g7EJBl+q1lXosPIsr5CyR22tjyHUpwjkyWVifL+/ZL+K
pgzIhoPWBDuQ5iqYhRKI3kze/Z8cLS4vdxX03+INJQpGw/9eqEm6rbGzvzUynvXBDqJN0oLs5tXW
9MR/0vG8jGW8RzsDlQOf7d+0BwOcIVK6bYcd5KYF4QepUg5UQ+UZWPh3uVMr0kKo+w+7MXI0nvYL
jYrT5KCpRpHBttHf5xUm1eomvggkhQ4muJKwO494LQfdhdXt1iMxt2iIhq1gOoCHHm9NQE/6STWa
5Y7VZ6xsPNeiPbfi29V7mAXmlsaiIya3HMUn9F8AlL3j4t7qB4t5EmgorUssBUGI2CRtA/6kcP/9
1v4zwaVHZdjuibSGfz5RmwyhOmhPyRi4q17CHhEoxLOG3TW2/voR8SOG/yThwuYfdR6IsCL+lviL
6mx8iHEFU0YlmSKYlAcIq1eSetTMBCIER0wOyP/bQz4X0mEQqKEpps3uYx+JDwib+7b2InPCdsek
cLMv1DQK3VvkEXHTRvldlMu+4gI3q74y2U5gl2eNX3Zo7HIXVDLqnLmyKS/AUkiIpF4lDxhg7o1z
RVm00GsSTWavnI3Gjx5TSynVPIWI2wYyO4dAkyVjWUaIyMHOy3fUicE4ppiU1CkxdYvo/WeENQeS
rwyauWGPZJ4rw1Gl3QgFtiIaBG+oPWAWJPuC/swkSJfMF1vO1XBkHj0bkRE1/M0mx7gl4q3k/gzQ
fLY/cHmsNmErn4HY33Ad6AXmxP3nwvuD08iLZ28VIFxkkOK3vmgGw0jpBML/yelQysXRIGKbCZzE
C9PjaN4ry3T2dFw/ZVUk00b9YGDNKWlJUX6w/5E9wIO38WS+jWsz5P8kFppOfo/Mcz+kjL+EvU1d
bIKtAEMgHjyoYMGzHzTg3TXP+cuJ3IyM0tO+S8RqwBDlhPLIsOd+utSOn0YvTWpbH8tnnV3nuLcQ
j8IK8k8FXjX92B3gTKyi/RGC/RpDy9HF+OEv0VlPb/DU8NVGcsWcuFLnXYASCbKwvQLNN7aVCjSa
3XyCVhzXhIOmrdmutLhRvEcp9CgI4BR3vOUHGObbhtyxnb/hVAQ9QEZeVTlAjus/8szvhe3t7ulw
xYoON7JDSAYVYsyBuNZFpjhxYkXmS+wDZcGHtr8fwCdUFivYuXlA7Ccn+Lb7RZmawAu3zm+Nzkbf
487VJ0SDDBE1noqPGSl14Wp9s2HMnApqAF44FgtyeN5IexMFsf9/PIQkKyWuAivAvYgjAANHbWGe
AHYN1z5zadW/f58u00eZiTnQ7aYAAB0RI5RMpTinS4LodhyPSq+Vm1sPCaUVEq7EUBptrJaVdDzn
QKhMW8JNGAkkIzC6sn8jgBNF270UEc7NnEKsDVzzYfJkiIjdCmV5i11I2TIAUv5Y0G7rIHXrSFx7
tab7RV+Nrhdn/g6Re+m4QweI2j7Dz2sRCUAWrmjIvyMXd1oAgJG9gJJLfg1vMXehltE5wA9LfF28
rK2nRkOyXlP5SrFklXAX6rbMm5iNNZO8DacxqtOJyk1XNAa1n68BEmNpra3+5L0fnx9XCiYut00V
U4BPUk6lbu9L4wbP4KYdyYI83IZGMGEpYuBsp+JiDLzWWuWc6BAenBUnZ5u7HDGmHt5npFFMF59w
zLUWAhXcVxD3zf7Jj2dc640oZKCg38fj34omhlj1KReZKLxxBB2Xp+7yHOS0cN9hY7ftOaRnJdO8
qDMSvJLVhpeqPWq3ZgdrQHnylCl7k2fCGp0UChBjPP4vspsNdXKWnGhLToe7nnGUPEB5wT1eQkfI
MQmoj6xH0LkkAQsu7urxXFUJI1xzzPO16l9f0Snl41ox01fHfrt3hZPQJMFTNFnEOu+F842Arblu
78F7SBGN0dUEocFnzFWR1cCSUlwVXpZ41U9k/GAqvalTlriD+4dUg1n8vUkXO66ln0OaBt9Q3mcm
x4dLkUuF/vvGY/3kyBILWpHY1xatnwzcJEGAnn0XjkeLJ+2BVI3jvKAa73JFw4dWIIncGKsEksHa
eD6TX+hMGWjIoFMSEw7YFtBJB2S0HrQs8N7HNqECpWbmU89jss/Hw0qvx4UJbABt08mOR3Yezfk+
8OGRoKw/qXY0r96B2rRzu55LyRkRqeIKn2Gl/sJ8trS/AMmIBfFCIvpWYxqbuVUzQxzePWJLSswJ
14EleORL/NDNKniXSHqsCkCtL4Nb+ezMhZZFBWxGez+SiCMLiXsbfqYkocptWOYTbPsy6LvfZ+nm
69y/Vb11d5UaY8kLcQzrgybYHNrS1YADcjaJorJH5YoOBICkxzkRNaNLXwZakeKwqL3EcTdRPvaw
aPfVCgyfmI8QT600w0/IF1D9Cc+KNGGkO7A2GJ0X59F4gjI5RNBApChOGVQ01FfS8FQXdajDTyTI
xmNyFkr6VwGXIbQmya5pPCQlAMZJ53Tud8gBm82gDotDsXZ9DiqLiGbyRsFvaL9qbw94ok7t91s+
e2wC27F5pF69fmCubnApIyCVvi+RF3VgFBGheOzLngJ1yL6C5lyI8aC6YhiTbfENJ8f3OzbmM0xu
CJTTTUEWrQRsc+eWZYLBXjFTKT9A5CX5v6mpHv7epyq9+RaIUD3dfhCTVWaoLotrqQv6hTZQh7rw
TIbNtTFDj4xFeTBvYVj6yBUGfXu3fP6A5V4l1XOB1n6/cb1oz1Bq9knWL0zIA/0OiWGisvW9u2Qz
oScIG//svz4HrqLGN2eii9CmEOL7epUuISnnIUJwi6vnRDJ631+VW/N2na1djLnXHrQfWUt8uKJS
CljXrjhprfK60saRJHt8my7LwsfsBVT4J/BZ5+AtnkrlserkzJauEMeansDUvuGtH3QUR5fERW5g
f6PeQW0OjgZfw9CbL8fscS+gUF9f0+OXhjnYWFhCKaAY9bJuPYpT9HkGdZdKJ/62HaMjV8ostzDN
ddU0rj3ekZEDaKrD0b+2P2sevYjXZM7j156LIBoiquzkchszL8MtDc6vUO1tCD/jref2GJyAQh6p
9bIuB3CYon9F9aGITMjAz9FYBRR6KcdJCo7wuRJWHI3ZpgjI4btzJcX1TT7gROFzcEq7Zlw+T16G
9AoE62FmK79rboLz6ikPW4hrEwp9Hbfuo1AWN7QnF7hxmW/lBX4hVHTAqAZL/khOzgmE0186fsG6
GQoFgik/+Pv1EKl+01GmpOCr++ApmSyE87/nRpu0vTK4wuY4KnIMJABa8rQ0PcqDqGm8nDdYXlMi
cvg7EatdIuNTVGpwN+pbgqFlZmgCQJkZfouWNF+gquNgziGcsFgv0UK8C6pJd4s/snOjZ1RnT2et
ZY9X+HVrVwrUKzMnjsCiXjGGTihavuc0+aFSg1f4tn7ZYLjpt04XYpCI3xs/zdoIB/qM+b9FByjc
XX0vWrPf7tw88VqVFme+Gcft7AzuuqrQ1PJkcj3bqZEzAM9I/jdCHoWOECY09m/WKU7Zy63CLSU2
jFsROEJPC6TdIJUSEdwqG+hzncYoXps0HO9eFNbkh1gW/SMMOFz8hzgyDeUDBA34ASTqAcy66UDU
q6P8DXbkxMIGqZHzrPw6GkXP31bAxsuHh47BwfmUbZmbgHtz8y/qtAIchyH9LPtyRTxDkSm10Ztf
NJTvSeuoO93Dp8GPOTOLyP1ANyJpy/IaFoTSVDrypZq03KLeiGu/28ngVG/QzElk5HBcvO7z/4QW
jsy2VWqF1YPw3X3D6JuSuvEhRfPeej731oPqgiYKJwm17G8XRRYVL7o9YDxElxIauhGwYzOdDIqj
LusW4X3gUR8/W70qqixfslzJKl7AzXQaTFoeNAlfKDpJJBVam+27bwP+yrbxwyXon/tfEnsLf7er
d/DeUdIb3JVKZCJgqjTUaAZeeXTc8ZUApz35Ze8exOfUMEYDUt2UQWSt6cofnsNjAyPYhvV/sXBY
rOoDgqzQhahjdwLyHgrRUWZj+4J3GChsTgIN7xpLV1Ts+R5O515LYkGhlHZRBwSqF+oAJw83300/
0NFFO/bXwyY9fg6NwmnnlxfTnvkPCz9rxG71zcIiynLo4jE6347PovGL/QlOgLThnCM6FXgREuy7
wptTqfW2tWi4GIstWX5g/36pvZTYmkWX4YwQhEnD227BODFzNM9z3GcNt8MfofqIS7/SNrN6Q5RR
+S6lRRg3reeDzx59xXIcV5/4b2xfsSmyf6j1hq+AXnR/zUkvEoZRKa0ncfl4TNvIG2l7S4nlBYjh
uP/mITxwSvAjVRA4UCLAyhtrlL9HobVAlj+wz0zGiNo9CQRUvKIZZ7Cj4k5tyQJves+REHO7kO7c
DFIdfBS/gKcZ4UA4/L9DXy+S1IHyGIBPBAsgXXimCi3n4BQCFcqSq6lp4vAIUODwr7E1sRv5et+Q
SpG8GauF5Q2dP2p5xxZU0EeZTv6xBDJ/RE560If3QdYEqyjmuisqiD1mJ+SkagQCj/gn91pgMSli
hiojtkZQgykoRxhwAJv3Dqwg7W3DHNKXbMwSqc68Mh3qH3rZzXYcXcMnDvs0FDOlNgCc53LzRtvY
xKPwRK7h5U4RmLM5BVC/HIvPPC9UMflXH6fjYNjDLT/Y8GA9eMNQwEJqhlS/x4cY7HvlzaLX2RUr
2DSCzmLBVj89naI1FAjxJofWaApimv6sIhzf3j4t90JQE7B4P1cx6P9lmc/NK8YWGW4Bqe70MgdC
aiiRgPnldeyOwYfMQDrZkx7IOQjXPttjJlBjtXWuduce5onByNDU4M81sZk+Psmr3y9Uol06Clqq
WkmetaIa1tyci3fJK2JJLXSdR6WKWrF4xanonTFibD9Ah306zQRbO6BNfbvgyYpCdLAsn1ORNl1S
Rq/0uiVe1ZTpjry1dm811C9vZmX2U0+tkHxbLoMrPKOJr7i/K9kqEcbRPbA+oZupq67mQHMYdj8W
eadgeEUzXEqtHAqNump9IYOxoj9NWfG9HNc9qEelBD5ORHxx4ydmCifF3Ya3lysoNYIHydOCfbun
+H68RxkuoDOKY4G5hJDzIHHTOloxqZD0YtK9hiUFayIHAOB9drX4019YnPUjq/MpXUUOwefX+Ote
OsRIgulIvMWlXMUHlE/s00goOz07lD/QlQwsQGhaErBMtPV877GSwd4rzGEuUuHoHNSnMz2IguXO
S533eBe5bfEAfPgn3RJTTGqTK8Mhhpc9zNWigujWX1YP1m05QkIaVq6k6tR06BsLjuYiTRyI2FJ/
h/AfQ37C1Rfc0yo53KawKiVpJhChM+/9SoJ+Bmd/KZ6z903cB16IPjujPELl15lHJJt48RE8TS5u
YtFfD9b+Yer+K1zCGX5Nag8EPvAysjjuaXzgiSWVnXYbUs2SJNz9cfN6/qGNeKuYVT6JuIpSXEB8
QYkdN7LdhvJC5PVP88ONAVC0FiAtblWVvvS+oVTikpweEAGl7NJ3wqlokMKZpjoyoq0WSIrDQnEE
sUq54Xfr/S/0C3hcStztYSp5SgFHYmFFINwBRN6Rw1BlEWRSR0389DhSICXk16wpvv/4cbkzY2bF
+Ivh+Dxs3xi0w8Kz9ab6d9DcsybxGj4SDuMEPU9lK1YBcgDkPQR1sfuUETvp5SA0b7nCon0Cfskz
WLOSC8bjjaoxyW/KSZLPROu28BMKQS81qvgF8Byw/FvPPzuY5gyA6MLg2QmD5DV09HS2SDBgm5u+
/Oxr9oezMIWmlqrX2YNg3g7IB7Y2LujUeiSWY0odg/ssYcMLSufNwgMOPZXia6acCP2xZUUACUhb
GVWC5UVjC8Gnc6tZm1242bYDM5V3qvE+dkZyodhfuXDaMOgnqTF/+oBgIsG4vE/ZJgSU22J4pcLk
HldCz/jLClzQzYbcEgL9gfdcFezX73+75+cb5Rd1ukN5fnliB0uEMnHN2Sflqf0ravtVMvsySvf+
GYKlpJDS7uPOFZWypwvxUWmPaGD6TMwFm9mccoKGc/LoMp3Pdj7ZZjOL/5qGdjTts/QydeQkPyIS
L1cLzvYpANExHzJK3+X2k7tOMoy8oNTvzwM3pZJJQy/opvB9DqV7ydsjj5cEbU8+DEYO7RHpxkpz
gygXi2NbnihGa/6ZDeFrJ9Z5Rc0KBLWRrGi1fiZve3TkedO0056UXAhpzWq1EsC0+7Y775gtFkng
WXvT0D5PhNBD3bqhCqyxhCSXD0NOG/T11YlevvwM5GvkKAB25Mplz5mYZZH4iWuJ7DysaVPSH/gB
gApw8gpGatzVBgDFt04oR8Z1rErcZgIVLxXCvCwU0rSjlaAlLtbHlsAKx7q+mfW01k3akQ0TPYSb
o7s3ZWaQyAlOA+emdgoMBb0Nzh9po0KToRp7j5WIGesa+KQ3clpKyWneDLEQWeTD7U4YxjBD5K4t
HoXIBQkvfPJwkLsTMRXsdo5JexYC9Q71K4/dCzlWXAFcCWV7jtc4oniUz2H1x0EwOAKuAVUFQ5Oc
yMV0lqJdazVdINtLQHQ/4/ZV6BxfjQ6de6NoO5rjwHcHli+3trHD0KwHIgNrESIcvHdaF1aJvdI/
D68Cmz0A/FX+DgcWUgMJPDbLoy0wQwT28hpZ9s3veJa44Gtd6ALQD7nNHVnrFUHXLi7O2jYW55Jf
+enKRrPgOoiuGHOreT3ToJcTUGqYEt2RtF+yRz8hBnT5YFQId/y8kZ1FsG59/1cPgqdFSOSxMjTH
GcQonO5qn0iHSMYUtQ1PLCsT5vEjkZ3iqPsPK2ggsCLa8Z4YWF80IwsR+1dWBRVukHcb2E3ZEjK4
BSYVwOTr3pPMe8OzPk82w6+0tFH3iT+pw8RlvfYPMyTthZHB8aOeuD96v7+Jf3fWY23WN/64gmxp
rq8178tCZ3S3PzX1cy6C5QkAnG4kadvW5SQLfl+SW6T4kgnzbe/+uqdGozogV+M7VoUtc3oSL2uU
G3hl3UHu5Gd4tQbcwrjIeCUr3W00ognjaMt8+7XIn6DHR5iHQfgqP3GTInDg6ABQhAIYXvr51aBE
U7C+Jq4iHf05AckmFohUoHFkZQ+F2EB91zmQ7FBIvvk08oZFwN9c4+7bJMYL0TkI0Lc5ZFC1QQpF
OzKGQTEBD/6tmYGAFLXZVQHeuad494dIfSa7Oz9xwuaWHW5dCTDWuG6eVjzU6UgsF4urQmP/C/FI
UPJUqUsdb8LHTsrryFBtxyDL6VSW5fiiKSEWcD4UjrCmwtiBkhmqCU5gElrQ5vm1egpEGExN11lj
88mjAF5gXTNcihct3rasz1Y3ciNHteWvQtpzmqeWfIjMuAlJdV1T/uN4bELVgG4TImkJCEW/jWle
16YbbwkFfYy2XqzIFIHaeHmezMiRMKIbGvLi7bODOCcIitErFXh2qQ9KvoJCTFvIlxiC1n48vY02
GaNIuHdUUZj8lsudPx37dlvt01i/saDmzuB7qLJoZSrpH/pMWlLAeshnwECu8kp45w1Cr3TwLCnn
/N5+XQekpzjxH4oo5K/KE/RlaZRFMm9do0FzA67i2o31vsKOdo4M3cLbEplEFA3ypu1oFnCDn5vD
/hSP2EbNmdht2zIT6e7li8SREIwuEzh7F50xi2FYYCiQKk3BDs898lWsE3HFn4gndm+wUwkaQNHn
dT3YiLe8DTXH5MqI2Qjpd5i5fxak3jHH1TdyQrXPenxla97RX1jQie4utRy6jeQ3ULWXeVP4hh7x
M3h/nRPFJ6WRJyXB1NulmIWAjChJzwvN6DaqOW5IyP8goqYYgplz6Os9pxfy6Y9VAUQFRWZmnu/u
+9IarlLsFkr3ycS1RXpi6NGSHkNaRNP4/48QV6ATJgAV7A8wM8CqTVamZyCBDuWQNzoRwfrUv365
ia/1TLoPLehRzZyTBzqdPLtdQ2x+KgsIuwOujVRloRJgsQgJym0aV3haAGdV5fO8nZKP7yZqZJpb
arjGAr9qqiBenKFVY3KPW2UKQGC8esiUX9TRs/0A6jeyi63m0/dBbz6ybyVaJPhreqvhHGujqSee
Cs9OJTp2fRJOYU9YAOXMMDwikIo/AFhq9PujcIlNXSgOsaCKnxOrXwBrcFSbUPxtbb3nkIJY2moo
vWcRXlKc4I758eVbe0TME093d8PZGYfQnFQwDcve/NKoke037Ahh4BLH5gwhxaRoCBhTGKHzwJ8/
Cpsfwsf7V8PcV2+/hkPXZMNcNxIHzKo1veJBHkwtXJHrYEUNOf9XG53urezNxNtijLFOgoeNtBwM
zMtlk9K61MbZWFg1R3ucKHjwu/DRY70pBiLe1ja/9M4I1QxxFZYoBczZOIL3ABk5kU8ElAknBTTB
w5f2nMlrv/miI9FSXaMfuSLbJCzVDS13j+aWWuaYX40tWS2ChNJwY1X4fc6IB4FabgglL/ZYfq2w
+5Iu8eENgKaMPTjAQYvynGXbs9CVC6usY8lgWXDyw0HRJv52ZqFsEgsfQkCiP6hkrxS7U1QF6NQI
8fA0q+wAd9+NDWTxCSeVTKEzf+QJoyXAAvPnMNbDjMwYJZIKnmcpEGNj46FrS0C9UlheIbjiP95H
dAGAoUd+XV6i7GXT4moatFJt7LMLhTw7purCU+bdnVSDPz/krN+sHNdEHix4ndi7G7GUx1XVl4PG
P4D3G6oKV8laWXGhokyM6dK7ktbt5XBuw1sHkNLdt/o6astArotjXdWg6lVXNFQbsWHuF701wyx4
Ogk9ds76lPs4U/h/NF0LscXldbgyAJ0Ozz13DeFrwvICq+HZoL8A8a+9EZ/L/YcbgPnIW/QAkLbL
fmBQrc5SqiihHJubAZ6QcfxO2mnBaTLuS+A+RD6NRWHEHWf0hcHRgCeWqp26J/4jswN/uFLTsKNh
Xc5EJMgLxtOpSBC+oBITV7SMmd7zNHbPyIqcLmXrGGZaf0XP9C4fVHIGk5tCQRw4J8v0ujSvOySc
TBPInVCQFw1y1GGSEQpobOFjbdZZy2btukjc11tCy+neVags02XW5FqYc7T0zhANFDaB4OOllUqn
y7/YOtCFbztpGjfSNc85Zf7HvMLQWM/6QuG36iaKoKdgYBmIyjdGOO/O4TNhL7/SHRtlTxgr9+sl
pNUm56RWxnoAGZ65tU6k/6zpvNgoArVmWPK2y9LZNKNE6zwdTyeCVYJeTI0VnGylWgw+QOTprgqa
Yn2aE4Q1QDsY02SMYYGWGdy1ajrqSQ2D2qR1EFN8W5xvyNVVr/azsC6ItvJ2VFoEXKJFeYNwMCJs
LWIv2Y2tOPYCK4M6y30hKIXixHV9bzr8jsEPZ0qPf+SkAqBoXrcEh7ixDyupl3VZ0q5Uqshfdxug
glIsStL5TwDJPnvib4SH4HSoGaJo20hzr7Y4FF6IUaKBqMxLRbQixiaGmb6VXTC/N7Mt0tFfPq+W
MhBoXMLkK1UV7XvDkvhB0GMiJeb63tYPVafNOjiTSlwEHnPie5ybW4z+WZtdMiWnpAJWVmO2/hIC
O955DasaMaG7qcRgejgYpUL+8Lu5M4rUip27cmrZe3ftOYTF/mxak+Kqpg+gX1JgyU2amr571xOp
bxBTOZalO8B4eUEbMKuv9Y1AbTH8uyC54+lfyOfR70ZUlZdb9tuLOA0FMo/AKh8gso6ZrZ0IVPtD
G06B4VS4CwXVOqN2iDayNokHflC3LNq+jlGz9rvFikHDJhDfCQ8Saz+GpuyKqMa7+xcPGCy74YQB
dAo+Ui56IjXQlblXSAeY66UmafNH1bgha73TdsbTw9aozFvfuBrnPb/XuXjOokoYcy3uhv+PW4zz
5JOwK9Xv/MLQl0T+/Gts8zjUxNKIA3JY6zRa42/M9799r1IyQhENSKiLb48k1B69zUxoOSP5+aqO
wLJdOFBBpG3gdyCS5Qv0ug3FZXKYUuzFIiNUO1MLLiu5blztkWup4wiXDBsMZzu3xu20wgw8I1XG
Qrhu0QDQtkUl61V//QGR+9Jwvq1SxRq4o/fmTHLjlSHTGKXqfGyMPwvm3dlekq+MlsDFyRgzj1In
v7+scZtNA8xxWbls43gqmj7trc0IMZEEUlIQQEwwAiH6GKxhSq4pdYj5wTE4Vso89q6Mu/V8ncfo
uUpHHE4Wq/9gsOKijlNCRe9wGiIw103P8zwHOUA8Wxpwc5Iptys7IFHKB+5fBH/ISOAFx0mXCeN+
QfskWsp8JetUUNPn5DGjNSUzqPss94RhQ+vA3KeETxmhVbYnSYyapc33y7tArsXL9Fe4nCe3rxe2
DiSnSzGGoPbSwTwfbqqXuht3o7hJgEOwKJii8XKzn+bWTHYkAXmoYJmxPlbzygQ6pNOfivX7ct5Y
ew4ZV75LHaQo7JN1uhCvpF+GcslwHzJzRP6IOntTQL3j6d2f+WDnXWvP1Hn8MNxZbdPTgcf/uSLD
tOunLGnbNHkCk2yZUbDxLyT5bRpZ5XSnH2i3lasirbEH7Gwv81vVWNkmlANKuDnqxuh6tYmt9yAZ
kjHuD7qLTBkKDT9tbL/1wherfsUIPLpC5wnJJ9mO1P4M8dpR2Qjp8juQdOsrTnoBWVBZ55Xj/gp0
mbYE+JtGmIFI2wLs1/83Zt9fXQGJjKnhAaxpMreP9Ovnv9qzXwbjPBqlUJ1bU8hGAt2CyrxwqXtr
OGsGDqwaGAE9QiV1BJTuFAq97BuFa/nagzH/tQ7cfjtG/UeINphq9WfanQhddw7A44JOAxpzG4km
KCUKNyTlFA2DF+cNJeaMOnYY3FqyRavM7NiAU2HcWgsYy/1zhT3vdKcSyjd1ZvuXSzcaE5Rl/lwN
FnWvgIent+RZY4X9uXUKzb0sAeng0NsdUBySGAY4ckXPYhLPl44mi20KKlwkV5Q22rnHabAKXXSk
6f5sG6tXwxttJUWflTyymgENVFweem0h8fjq03lwRWJigDJZdRbhrhbnnnsPiMsxevqb1X3EtDvm
Mh8Hq0DWhOvH/s41ej3KtnJcOn5pu85EKno5TOX+hg8RpgXPXqtlhvAxClcies4VMlEZsfVIKiJE
Q0rChVjMVW+zrKHwk4/b1Y13FhbCvmGGnL6kMOcFkYHhNEopD5dkZzsUJq24jk3BdF6q6lnewW6Y
kLuzc86eplV4vA420o5xZhvd9B5eoA11yltpBIuR3ubVJiF1oNWmtDHiTJNdK2jc/dtO6JgyF7pE
29v/RcQLHY6083DENgbFP8+QUIruoAb8VgJlSfdwfgSatnth3/5aQYxZ2RW6eUX0uiBHFZsiObPM
Va8WMkF1H8nntciSiv/4wC4i2K7IDK+SqDeFk62ZiGvMWO0ltaFxqEGGaGzs4MHdizGxOM2ARVq5
5MPER6NqhmzWfGVKIInCzaLn+IuOf2KdPUAdUnHL4OBQJLZ/ksPQe0ZYyxIofFHohSGSUEneh3is
PtLBf8fHzB5m4Dm91paXjfib4noPPHZ+YOwfpASDUQOZUOZUc+wB3jiIrr/sGlEbKx9WcBvMkMWA
uzOQqJ3bTOpaYSplI7dE+7YQG56yToG86IFuSOoCdEQ70nTvdc3BbSCHr176yVExCVu0PjAQwRhV
9uzH6n23wo5hGT2C/wFLwAF2Ru2F4nNYfkNrsDqrhWFznEwmxUsvPYj1CdFMD390aO00hwuzsCOJ
PDmucAEB0xpAOEgOFfDXLdamelSONKpD1396BQkr7tJv7XYApG1JgzaGQUkOjylN+YBcXy+hX8gA
39biBqkiUxcViH+w0d+DTEPoWEPDzjYuxHZvdBSv/an325eQNl8smOsWDABZ7g8BxB6yMsXZZVNM
ntNeerpk3GyVriPH8UW3NyGO86wFi/p//TTV8J4f09uYez5Rv1i2EmyaSL60Hxj2Z9lZcK+RK2mL
R8oq+G9ozFyUTrVb3A5rbuV8KIlGYRHfz7g/z3f7rG5jDQn8qFiDEnDTqrWTMfx8CXD4EzAHK6VW
5bShyS7oBKjxDnGaepJfZAUtjy0pcspSfrP1eeney7jnGbpcOJC+5V2Ds+mktWT+lpkEts8dyf7K
90zCxYF5KHV9xHSpPlfEL1wZUV25XH/KzY+wfAL9MM2ygq9pJHPN2TnA+Nmgex0Ki5ieMlP4P2II
kKldNzmuaTGdG99r+hZ4incvvulBUFof3BHjG/6e8FkPdWaLyQsXybeWZea1z8+6K/VsC1LNNx1x
BcV0qPKBPabCkXDcoNtT87BDMX5p8X2Vx8WACsAaqIji9uYaCrEwztSZqs+TyrGvPQFnOeDNiE3w
D/Ycs3GM4yJhBxOwgafZWMkXERw66HIuvbvNXIItPB25kmqMI2UpNl/b9UMKzVhg/fw5Q2jHb+yv
nkis2dtZGlUlhK06T2Wdyv5rlAGzBhSzG6p7nPMBysYlBOuyNve+0hxzBNwZl1UUxxhzQui/JiZX
1rj2ja+S5erRKYfkNv8KeDl+Yd6ooA5+ckM68GbGMAxe+T0tcq959wUiGQkKmIgwDcAXoZA5gOVb
fo50x0IWa0TDfjdBK/nS7TbigC6ee8+FTXPM5wjNpMAGcrB9g0IaBHBpKt+GNPv6MB1zhMqaMbW9
Q33Ncn7t/VrvohNreD/tPRf7jxPZV6d3Q7hNk54+dGWZUWyjeGs//YAgOYzpPsI39ojVPrHIsJkz
LyNZL8yvLWtHf5SVZO5tTa/Gg0KUtAuYvKdCHfB3sGF7Ov44wmViQiaYzfuLzt7TbXY3YGFgvYAe
RTfcTT/Z1KmIrkKHFrXYurudVj1rVk/lIuzDR60b6QFtp84r8h+QMhL8CAdkNJyeuLDaMyVr1Env
Tjsqpmv/ou/PUa8uYYJ76KB7DfhrmwQ7UEh6L1cRsfNadTh4A29vtCoO7+hbWm9L+XPBFNIlmadf
TDlDMVb4b2+2awd2X6kz2PvNF901f+KxpixdC7owIi5NYEI04vqCtJ3++XCwvCLl55Cd20WQvYlR
mcVSzwTS3JuERkpxpHPktzBm5JVof83YeUae5mI0qjgopt5fCFkkWiPIQdCrN3y5uDmpcMc2vDpD
aoE4YMtvBZfc3X+OswzTA/C2jaM06GMTNwzomFbLhGvkpCtJmdEdqupDVdw7C4tM7uRZODp+9kln
wigmoCfTJRhgMgRq62SiV/3UbbImlWYJEWhpkeRB9FEk+rP2exMvlADW92yPfOqY54LOJlXHqF4h
6HnX+R+IIfD6/ygrOdwCZifSIRGf10gxu3qqAWX4cygU2bEVDLDggYQN6qKXq8vuRXtA2sRYEhpj
y5jFXKWA+mKjjMybYSvwXAzuDlN4VYmy9pjVkUkVoJ3RvfxkD22ciC5IbYWXIT7sF28WxSFCIfOr
Jl7D4I+y+9oTMnXjxpHBwf7NIal+yu20xO00nxcTcMVM5wg4gB9pZTs9WgQEw4zWmbjwynK7wsSL
qTvpXj6tun4khIdPzqJ0+JEiVu/wBxG5D7Oi5VdiVpvoU9MwW1C1KpgaffVg3FmNsd5+hJetVWDl
PU+XSxcxTWPIts1loTphSZvTree7OmZ5RN5iOvWn/pT6xt3lEuxHq308DYDosxo//E7Uw3YB67id
f7MQ2yiS0K1YE0ypjjRQIeQknzwi+dlAe89DMZXejJZ3KS9TiwMv0hkaq1NtmRfZ5Mhb4XUScJFX
bdwdUAibxCJqabpsdbzju/0341sToR/JwnHmlztc1R6Sqsy4WgMmfBn2a7mhI7jpUAksz/iQ4QPI
zOLA4ND4hRvUs6xHw6zaheyFme1VrDI+UzCzvB5+bx6ZZrjA/r7b7IqpYZkoEvwrpoED0OYoY8s5
9HjZ2TB2FcsaziUCfWLtkUhpAFYXu3n4JqI33z9yxfhwY+ZSwe0RoitDiT7L+S+IVqwHTO8u6OK6
+vZrvSaZ2lk2L18k3pklYAXhpXkCh0d1mvSGsHn57fBVbDE9zHvX1O9ba0TdUKWbgXA/Z6GEIJPD
fAQBg7MDmPE3LGpF+QcDJ44awiwPli2znhmv6kBl74Gr0/AO+1UnKHHcl9TMNDfVcUPqjVD4jdBM
YL8p18j9dUYOq7kiRWr8t+8J/VOMzLL1ul3ksN3/gOi92or9YjLXUl7qEj567hnVC3P7chJS9fZ2
6K5bTitLOZu6oZmXAMAumlbjjTc8SUXhNgBDKh/nQpMItWvrlO+rO4XQ/GTMmqPtajYYBvhmL64v
ctj0BCA+T7S8wI+xF4KI14LEA6PFe3yLhh9fxW3L2nsrQImZAdB6sKca5F9mvKbM0UygopJdbSMT
cWOxcgtwxMhDm54eTtdbO3rKLhA0JkRTmUy9zX4yYJCOjlDRi6jkKKvgxSEXAdOfMbjdqLXeHEwH
yagUvGVPGYM4fVirhWFK3micGRpOXyPyy/l48Ucoc/V69OAy1nf5UvtqmTOiul0PMzPnCx4xw/dp
STPoTRzGTBoUf/rARZ/c+7ncdRn5pqC+kSnQ1/qZKaQQ6CwxXK9w3iPEQcTXoa36Dsh0iPR2fn6E
zpg0LexwUi3Q6ZKRooQpnuFdy4/Me+7YlbnZ002qRP+P227+JB6KKqce5Hu+MryiOqGyYark+/l8
XMVK0L8ztnWCbYP9VePh39e/w4pjM3pRDCO/lqZ0Nx++cvyNA2o+9OAXgwHt/lD+E2fbFHaUpJ9A
ObiTU5J3yXJHf6mBE+zVg1omF2t/axyvrmJVC/t5veP7kQF5vM1nJR7JOK8DbFPksDuC7D2Pl4Uv
ri2sZXKalBtEmmJK8JE3/GAb4IAQc9nUTvVCTZyFLtUKehXtKPk1X5PQYRrdxIVkQlcOeXCCBrTK
4EzxFGAbwtKS9+9vLpYDDqF/dQl5gcum+pdArmoGQyhU3OrPi6mgi0whZFJXMomJ5degiOP6G/ke
284nvcMH7ggxBICd2xHcWaSjPUQofuR/OX4BpTVO52xBH8EgM3w517+fL3MW1/ZYDFSyx4X6X+Vd
Dh4wibaXIgAMDwJ6U/piYcpHaBQJuGcaQmg6EJjWVzl0vgFEPL/bpVQPfw7FFWXMMEdrU5lNek7C
QJT3WOabRA1C3Bv9h126scGG7Jnv0ilLLUa+yZWxio5fxdgP3uh7ash4TeTahIWs7rea2IZteBHc
8MG3rQbLqWyiNffurjL2dc5xLvuUk+V79svjp1th7v/XqHCY3XHQzDOrS3+x2uD9TpvgDHOnUrKZ
PNeZD6B3xeGTxDt3VZJqo1Ja0Vf5BXPnoCgR2BV75D39SMhO1q3wbGN69eM7qBefS68GKUhn/7XF
qfLxw2kjSJOdWibMGfYHfdbCBgVpa5flYmIuU0I49YgAxIRpqhpMvIOUIqUCT2yWpgtLBcDCVTCv
WuDf6TLx37oc/5LsbUZwG8gDml2PJFrUkksSiuzON7bPnL0vidHQMC1TJGaTR7NGSxZ6+cGgr5Pg
dvrvz4ZLIfHkU4zdojkUv4HppbW/ScWx/UPALm5X8zGQHGQz3R8UjWHWTrUK8RO23h0sNvHp2nha
zH1ki8G4g3Vipv6kpy5F6eWTuMt0ZwWvA9dDzC4W2gzYRAd1AEtVyYK+CGEmFFScgAr8NiYkuw3u
JvzRxUSXnVyHWW0Mt1IfskEBcJsyTVztGWHlF1ppf/zsn9oLn1lp57c5SVAx0lI2Tu9vEWvc7dRr
HBHrGRaeuLmL3Xl+qda6B0IfN3+03uKTHzevmFUcFj/AUoW4W9LHQ8CA8OfmCycrdur6kWFAhiUg
ujkCMLs+Za6xIyauA2RXa046VntMkh/xXjesXbfl8i69IdAefnohOF/bH9DCIIQQAYF4IXv5WHlN
kEDpYQyn4kf6joBkU4pwkP15npf6P1dKrm5pI7bk7Vt5uRbnwT0BfLy5IS8WHRfXCzM2Hb1S8MA/
zJGjDeUk9lA1rGJMz4eblHgUw4n4DrkroHUSeCzLt9oCok2Vgbza1WiTyA1H23kd7flusOHfSpTe
MZV/sOs2ctsXUJLBZ+D4wTDoMyumot0Eo9Qe8kzLEQaid01mVL70lNVlxtHdwd7jBSJReABPuDnN
B5T1BprIR2eDHfcySf37hvij4MUV+9viJPrgJ4O97FpxTZcgus6RUjThg8yPhT2gurOh3pDdKm/f
6Ofb5s6EeUOG/WwXBmAqAiwNioGgKczNy//oVp+wDtGnFio7PsvYMGcLXPa1ciVITYCJIgFBUlKE
IRGT9IyHhyBOQ4F4an0Ut47oPzgbPUUYzyKiN4JnmZ0fQkZuxTpBCG1xs5ehBgUGY3to2KVBRXHs
prxGB45kAksTRbGPL1/myvxL1dyExf+Np22H6vaS4CNFgPxxMYfBLWTptszgbale+d031uTNh46D
vNbDXMA7BUZKwecty79FJ2PiK/2MDzC2RAI4njkf/4+BqIjdCYg6dDQ0/2JangiC+6cabtkQno1D
U0LtfEzA+nNIreodz2tR6kBN9lf+W8y8RuPE3Mp0ZvtB2lIzM3+LomslXV4InNJd/a3Ur/y6XUx0
o4RhVONAHn8PvhncHM0yC/IuFHPvCnU1IsAs3bkLMimepe6ljz7tD7J4nfpwiySzz+GV7rXB5VAR
u2XjV2g6pDgeKW5pwvLkatkgQfQY1CS5wq2weRDYRmAFNIz8DDiwQTLR9Q0LU0QYkVvYAXyN+sbK
uYsiZIbheSOoSjjVy5PELhQ/Hjz/khbUv9EhE5TH3vH+HMaekcOO4JDoy6JscRb9L/sc1ZEBgX51
V1fhwysT/giNKhwDxh79/1TQGnQxP7DRrK5WsXZvm6qTGE9OQoN3SsSR4D0MF8FCGHUR09HpHElS
6ueJ4fk/4ieG5pb+hXYgzrihrAcy3pnIU9yq/MDg7ujHrrRE5e+28jdIAxfT0R9k6hJrzv71QMta
kOQTAR0r7JygzfDeF6/skTT04xhGq9r6ThuzRTY0+A3N/XXuLADX568PlmaSm6UEs3e2ZU7ebKWC
vor8ThdYbBcdUs8Ae4NrSFwW38ictrSxZNOgRsjzm33fhaOW9NBYaXtugjBl7NhjDbDnJalJdZyV
hqeeB+jRiRhOYAalvRc2QgU4MJjCV2Iw7J+B6tdR6ozC9QuPu9VmP5fb0+OBoqeHMcr3e6cAn4iU
Omn1UDu1DdC/wHjvmbZa4BobjvjO/NxfgCPAWbBpTW9LUnYzRaMFwWB1N3xGld7gxypStfjCzqYk
KqfYKE9djqdOpVh17wv58BNRBpHYbQ0aRPtQyBGuWnD/vEhcdTph+iVtxdn+WYH1KeYpcz6B7RhO
QWHF3PymnhUVVRzUz4NRKL8XmNIjbccp0H/hBB+hyjLP8QJPPQZT/kyGXGTWfCPl1zlnM325kADi
KQJq954m7wzsVWtRc/cu6lIP8ZoZYvARB0LlNBfq/sGemrdL+4zX5faUHgT0SN19YAQWNpBQ7gOn
2UBOKf6Gv0vZTN1IoE6329rvUCuyPo7CSvndyim4l9J9tOhzeUD6YrKE+VyEzoAC9bB0B/ZLBElx
g8p68zImvqI+dRj6f26TdXRlmEnDZ2Wv8kq2xD2wa7Wmq/Uxg3IrCiVqY9MUapCj6d9zWaWQBU4m
6SZWL6o+5osIPpwvavMKBqqqMIfXML5KohhP+TpnZ00Z6RwLa/23/Nd3Dp/I3MTY7lZkd+Xvk9Rx
jCuHGNrvJPTXM42F7XK5wyQ8YRm8ynfuwTbtGSbHuj6MrHjqdPlkxY1AfJNjaKqYYt32UYGFK0Ur
1LtF4/9U5kddTunEqh0ZDJbwm5GDvg3Jf41x4Kzsj+84ioNC/BfIl8Nf9ap3AznA76zrT4vOjwq8
OzDkMp+KRARnZiurPslkB8RuHkwF1o3WeQ4tcNza7CRSalkM738TWU8Wme53FZJQ5c1AL7yXtc58
Vs2Kj1Hd48TJPR8h2cf5IEYuei2vThtlD0OKBz8NM7nc2lpMMuSLOvLv3q6bIz2nwatNt85FZlg8
uIHNfSgn7DaKu79HKRpDrKGn+0Axg27lSNxHxBZEwqHIJVgOKziof4qWyAcyWRMH9BRhmVLLLPsr
S+cO4r/28S4s9HJ1ogFq0X2CpPN/dbVxKNiOSf9UpX7i827VT8LlmzpFIHE5urrR3tBEj/zA1GGX
SQNBNsGyn87g4oSvyMfAdlZh1Tn2/EaKf1naNfxjusdEUlVwbT3NcWIe4vmiK21gZe2MEkwjCLFt
WwyqMVahmTrdZW3ntz7K+d6qGhuyVYWJeELhcvoNmzoQfM9ZLvlPmqZQpjnvbuE3wW5FOK+bUwUr
wVSgOa9VT+vHzw9dncIFGB8JAVcguuMTUiCZZelhVvzQX4PNiUkPNF3NitWB29uaJo97mYrx006o
pgNKydvkebIbvPNjMBITI8dxAyFQrZXnWKCu0EMNBdk8aJg8W+pYgVfD9Y9TVAf8Mrt1qMlo1uYU
E+NY5IKjpBOpUHmT+Vqr5WKzoTBgu6UrtY5FB1huu/9pVz/3KYOOhz/2JQ3ePfLElTBD8P3x7l1g
S/OjSj2iBFGJsm8E1ngLZ9j9jd9TuzZcA5FB6Ja2ZvjO+ZBEKr3CGnRSdznbjEUUNG8NFqjXnr0a
yJnK1XeS1XhT/TeQ4ByvZaI2dcoIdcBl38N8VuCR8hYKt03kzrrKVF88y5O0NL5LaaogSOIKiY12
A6CpuG3zVGjhhn74NtVXF+Ho7cBiB8M52jhlM+On0ga4q29j33nzSrcPQT1y29OjIDTTG+cOkrXF
oh2iLGABtMNfCUUA7C5u/kOnpdeujHRs2Feaisw7GIRuVVwfo9J4VDl/p10i5q6WFzB+nctyBI8G
DOt/WYLd4sRRUpAZV6jVSLODg3sGygTMXI2eP0njErRmbUa4gQEGyJfXVDpt0Gnkb8HJGtMwQ/aM
eaTPzmEpWrbnI9F8FLInGbNc/HzGwidfBMdHdCYvZLzr/W3tVFhzgWyZmZnNcYxh/7g4Kub7C8wU
qdHYibIURsIfTRoSEdaHs1yd331so4x9mPYvS/Y8QcopiykUzAnkXPdudYTC27VlYlwMGbiVRl2B
hNFSr1u4f3QUH2xsrDPfgbMUnxo5TcPQv2zX2BsgGEp93tnxNySSDOfQcWadcFhnRmDXgAmX+KYU
lrA7mCKxFyi9NLJs+E26gheEi0Kr5MToxjBG/wdiMjkZ9efRJLMahDtawxLU56UkcjFAZM3FsvPP
kRLV017uV4nGyB+PAhcZhu6q9xhme48A/YVp0Aje4sghx0lVCHnCw/nb3OudNb42in3TjwbHrkvL
ZkIXNDqUzQSXJRPfbBbXBqxqJhU+HDS0lWqP3TK/yVVZMCeVmIxl4sukR8GDfnt2XfUoKCf1fnn1
d7/lKU/0XdnZ485CEOgzAnVte84bykGrRLDxJWirfFmealBkjBCAd6FuVFuCslXkUyd9IXkJxRxk
8eEWSDqKcQSZ2j9Ja7GIzIEeU+kCD+Hu46qGt1U+YJYcyFybWZ52wEagPZItMvmSBe9u43lpJS60
IcQf9F8SlYk+pHq8h6fWrJlXTpWmLdu4ljp3FDgmlF++8OCbOVKdRrLjo8jLgwtCF9ruIqAZWS5Y
ECzg0frn5pafsH+IMQkKUPqjPKL7cXLKWwIrDlx05NXIpIKpe4Uh5ISq3WDPbpcFEteEmd+h2zxh
2WwcmJoujhnvpse3ovvSVQVidcYs0xs7U7uwZgtU+Z2WTM8LZx4xOdBqfdnLvyHRJfXi1gsgICYE
2HDS92px6bj4VXhVCWGbY3J29FrqibsAHDERidpcKpRERWa8aQEknVydvxnLaIUAh6bgwRSoy0Lp
PVRZoSGz3m7WYJD/jjLwwToZ/R5+hqwgZFAvLYSPWBP5pt0yYYPMnPRktaJWX+oo0D2CyWC0UjR4
ElYxltr3vT0AQra9ktijlz1I3r50uVtw8pnEDrpnzjznP6Irrk4iCzw9HL8xK4bTw9pr3jIlxl6w
qbXO6XMroz3fhI/BClz2fys1Bmg6a1H/R3MeaIqjHp9znHoc8w7D2LIhNDfCpAIAtJ3mCcPcLMbp
iYqlaPBe/X9AbK8aawh+QQCRpQN7YLjBQbPRLgRPT5S0mBuLTBQjTccLui8EJbzYVrk0Py2S/bUw
wN3WAa2952sEKFkvr8pu+dMtg9rhOFNG2/JekLd3pqA0nkNMu01/72vWu/bB2uGUtv8VoffzGEbt
0wwsATmQ+bWIxUZKK6tNdIHUK8n/M3yf80TSPj+yOl8BNlkJ/hwgowJlXH7YAtJL35/7vuxzawUZ
nEc09y2SE1bDAIPToq6cDragnUmpI5U8DjlRx5xZ2Q1E/RAWFqjLypb2/F9oN/JO5z+PMvTddloz
rkSGxR8HtQS0KcQMvLHVv5LwoM60LXnIjsW016NWu7diszBv0nIDq366OUNf+r4g1mv3gg1qq2YX
zRgdOO3X0zDP09lJlyUjrgZ+zPncYFs7YND0VLNzo1p6YleIY95bpNJJrZvsE3JGKwqdbYZgSSyK
zLY3ri/cODkmlfkRNBYkzMmsrvxJi4toGRtYeOAQi62p8BFTWleuqen7XB86kR+DSF1zG8996Muc
klwlA2lAjm0hLyUjsVbW6QJNY70VQldH4GyRR0E3D84mIYIIMgRSfq6igF1ZyCJtq0ZDG7bTeRxm
UKyZ7XNm0M0J1iiMS7R+peFILqukvn1dO2QKkhm9AvzHV1GsXvzOzZYRezg33jdmI0aG0V/8HOsP
bJby90zDKCRkC6cS0j5bJ10kEqVK3unlpUuN619MwAtRHkx6/+NDQr0RVg3Hg8qQsiwSj3x/LHqq
+aZGoj6jgkDJFLjWRsSXoyWSGvMoWuXjckua/S7L5rOBCRC2CQtoisJsoy32Md+IE90oOdBw0Rp2
04LxPD6zBnxWZOkkeJ+GpE5sppR/YY90Q1oZqwlvWK5Wmxfmr6ZlaZ0JrQneAUvz1bdcSMsxLdJi
Rt3uYe8eeb7wCq/Yk2Oiuz6q4ksCW1qfc+t0Bj7Nn1LIurVBS2wl7PmJxPCOQRcTRxeNL9/8PnKC
ELthiTk9opeVtLRrfXZRb6kX1FBEqFUQDuCM2g/McU4xuL5Mryj3x7Bf1XtdTGLYkzSDgn3MfyYV
CzSTvfmQB1pl4WpMy2t90s1vr7/V+HARXVWwaXE/qniIjQWLg/0/d+VeB5cVIhVmRvIbPcnuph3g
E4Htj4FokfWYCPU64ajCaPXx5+7pphtBh69rdWay+k+Scrv5wU8ZJvRkOoWRZqBdmZC4o50R+jCF
OFWRbcEoBUcX4Gi9C4cebyv5zRs7ObFL5fHbx2pVSfwXuWwET0rKhw/sSsK4ADt1NGFegiPctD+N
nJTy/DbLc9H8njQBZcc9K1qk9ai+kpPwFxcl9rY+o4f09ZVaU69Eaa3YsJ8n/gOCZq6qaIUrk8NO
Pa+c7IeiS7qA/QLTc3m/zS+Co2B0pcmvoHEGxvkKx6wmoP105jCu+8mlmUi5eEwSLPWi9gfcVN5i
9RqMcZglPSfIxgoI6OPYmVqhwrMMF+8lvgmE3MKwGSnFbiMMbYbkRzzq9YTiZZV9b+JimcUq6R+U
v1IButqxQgCBsr22y1TVTen8EKpjlQAGr5GOH6l7HUoLm1OpxwzJ+83NYXrRpB8sB8jiVz7BJbhy
4Na21HwaXwA+Dn3grOsvi24gURrvn0NgHFV7hiAY3EGBuLwWgkxiPvC313tEqIGarpTvinrsW14E
q4d0sp6Q1425jHBsfVBID0YLKv62WM2iGdrvgIJjnXb1rFHOYqb7nh9yHFNhI02G1Df9mQxkM+2/
kqRvVphE1A9VB+Hoo5NkNB1GYGm4YF+Deu0ESUVC/lqVbWJYmqJIO/FVwiMhvUXVonL2mQgHbXz3
pNgYri+u71gw8jU0fm/D/DkFPX3llQZG9HnEFx1yaAke1vscpfLBsy9apQNMLlahBvpRCpyPDtoD
8/0lvwA1x6GV1g2GV6wnuWpz4sBAUEio4i+NXSH1uJY/y/pV6Ue6616//4UY1YFHv9T3uT97Q+H7
M4ZX6N6NRq8JH02jfv1SULzbhRlAM2GE2A0CriW9FFy7QEdpIY4M52R4TPPLO3FAJeP7mEPifop7
ntuMQouw2WLKZBb7RXkywHV4ML5SVrrbgfbKSzbdH89GdZsirEKVIbQxU/hSUIIZx1Ag+UOek3VZ
E2y9nhjN4AjfrGpcGDTu6zau8OXo3MK3J2dPSs1U5Ip0VLXcuMhhKm73ckhZBqegxbufMB7QQWt2
3MfPy8Q55zVp5GOIaViNZpHcdnXft0parFkgCrJzlQwmwqKV4uVsZzouU2m3ddAw/qps4RrOkiaS
GcR4kbz+wW7HAtpyH77kWrqOulb/DpxRzwChIYTOswpy/35JWWP2LX8t6BKbjISRGs4EurapB5nX
FfDkhLhw30ApSpN0sn8JkiHggroXKwrAk8UzAbZkKncdEP1erkE0/41Gwtye8qkaR5QN0oSDF75j
xVjsdoL+NWehOYvGm6qzeTfTmSbS5+8MR+eytZWzutFt3deV/JM7fqN8RWvfX6uDqo/+Pz2W84vI
lMW4kRfiijf3SmnHe+MkXmqzarrsWn934xcc2u0tqgzvMM1A/GgKGCXT2/ZjE8GGAcyOz4vYUNsw
1i6hPEE9wVdPllORJwXw9cwJ5BcIVqK7bE+4BTmqf5krMBJMMdhgfMqaB/d0JwDl04ajcitiIr9U
O/P3JJk3b/ph5Yeemsw00HNXwYUxlP/4Buou888nzDxkW/d71wxcGPoVAeD9bxSYyAOvp+FKOrKZ
L5aVhe68R9UboDkYtlp0Ci+nq+hFRW+G8gHGLoKVUo+Bv77iU/FJPYEzRD7whmZA0pVVhaMTwfOW
E2ZOaQKsSH+iqJZFp1pWhNbNoyYsIYjfbuuZg1KPGTRxR0xpLfdpfR6pnwxHIY8y2iAfZ5WYNU00
WqVuoagsbbuDTHFylc9wKpdaoOie8vKf71mKLBGunDzCA+1K/y9lmqDkE03YD2hsFnoO+pusp/os
S1eRO4gUNukdQiY/8gSeX6EiHP+2ymODgqSLPJt3rxK4h/pq7AVpWmeBJPu1W7me5RMKDYFBD1Yu
LNj3KlEc77yCBIHdx6ZQ/KZtIqIifC8SA+fxDNBorRIExc/aZwFmyQYoil2jwoJsUDAr9hnoRHvL
FyoR9QtG3jnDMTgxY0CO8pplsWd6y+9UG8RIVJtxqes+PK0tWhJVKTRn7JoZK1tn38Go5l/cZ1TE
xYTkhOT4nRtCI0NEzDvdq4nqHJiwbt1TDPNANyCpb/ZMGg6DTde606k/njazPltQ7w0O0fOPnlqx
pMv9V96+Xx659hMfaurU5J4wxtQ4LxbgOxRk7xsF0YpZkFX9cZt5Yvi8iMvNvfkjXgB50h5ls5eC
hDCpnmEoEk8Jjp+GHRoCnnoOOFC6+6PW9qY0T5Ptwd/P2a40JQxts7Y8V4ZXv/AC2gmv8lZoMuLh
KWAiFRcb0vRST0I5UiH9jnuYjmw71FEgGCC0ztfjHbmElMLd6zO/8SQzCFhv9cWef0ZTX899E3fi
Hu28z2C3/n3gKkaVp54P97+i8Yq7I6mpgqd2ym83RbQgHcNGOqRi9AG4cP7eVaB0ZrgeVQRuxQGv
X1XCo/qcJHowx7m3anjVDKjJbndFvO44xiEggLLP6Sqxon4vxnCNyzbq5rX2O1nfdIg5XNWgCQKh
fJll/mIWc+Jp3BydJ28Xy7bH/gnfXz8O5w3KOYEdmrNveEzeC6+cDKtHOuamP+s0224f8cm8i8Ri
o6Ge2eRkJaUi3CD5QKKsGNYaaf+PYAxRq4yrE/UYgO+OGECj4MLoRL9b4doulINSNvIUuAxRn5I6
CbLY887+YmtXQLChr9zqVptE+YmN2Uw05UrFVJkBcaZgLTaH3XZuXEBx+dxnL7LLTNFX2uVVpsQv
9rx64kdU6AFaJHDqQxKjbrEeRyTB+tbLy96NsOGBQa8dEQyPZEXQeXs1fM+AKpKt/SheH7ZVIHeE
icZ7GNNovPd/XPZJ98rhVb3UfE8Ws8OnGGM+U473Rc/gUacni+t8qJHgtlf0ifcQeGu/5B/3FbkM
QTfdqlslgNWT4Mq3IpmIFAvVBTDiWLXmzDuSwDLdehKFtQGvUz80FeoGi3q/ebmtnyavi7/+lo+z
TYeq2MhD0Q1g4AyRessD1irCbMrJvx28rAL0QFZGsf7iJQ+T4hvJM1k9+G5iQu7n5caNq7os8QCf
u8QGkEIc0DIOS6/7LFtcWSrXEyIb29ijoU9mOE47EYO131aoaMKiKzA2eijTT7aTq/KBpua0yDnT
KVl4p+SCCiGHe99v62SybCuw4fL8X4Hn912Djy0vfJS9EKIqf2CtHh4jhktari811PWCUP6cx1f+
VyB6ubp9/F4hQBfAg1kBQcWFTODA5U2nmNvjcPdZab3BN+yPk/om0puCkfWyynpxYlGRYjGS9PIZ
Ne5djsDAEkAy7dYvhXDAOV5Zo7TYOfr3TESymrjCPjy8AyFqYvNNDfbcZm0Q80lNvzEfczL15rSD
es6+ypv15mdsQlz4V5KpkCOaRg/pN/lwW7LDmCFiwhcqnDHOKY+ELlNaQ11fLCnBOkDHgcZqmGw9
yUujGVAw+99MXm5pOismQnlC/72K4bQ7/1FyMGX52QkarGHJagyYRgyJy2obaI7h0luLDN2p4QDB
/Q2XcCptZWdfinwwzRS+Zoil97DXBNWDp53LQ9hrLxb1IVF3beFQ2pvd00zzXuFdHO//HZn0t/Ln
CPjidX8aOm1bdJ3WLeQqZFC1YXZiEvmd349RFMgM98hHze5rQ06I54m0JZd8SltjVlOgQwrw7Wa2
kC3yu7cFQUfC0YGOnXdMlhvNSyI9BEISTdvfovxRbYMTK9EqvscJvAZP8jgWOzOXevgR+/D1uz0H
QYQ2tPGTQmFMRjBgNR9fqIX8vPLFrDHPGS5b0Te1tzjgzMDWQPfcp0IwqX3c2w3NwaMQ06Lq/KC7
u5VEqD606uKJ6Xeblxp+BaP2cERvxBwzvxjYuBi3cGbo+e+dJRyeiuNhdYa0ChSfUxsW/PBe+E7+
HODEEKWfha/0abnEZfnucq+EtjkYoF76gseIVDo5sinVoWAFF8o20La7wRKUjfB8HGRlDLXjk6kX
2uCkO/bd2M9ZBEssK2c0DtyE4IYTJ7uL2hxtyrqd58jekEDjvBCtpMwuzrFaapQX5OAEDwXZ5CJN
VO0/BySzDUlSBlhDyQLrAEmenZjLHjso0EAiR86KLn+FUb5JvFNz5TLZbuijkco5nPQWwA+inZFx
McjfPW4+kvzBgp7k/Wmy/Pwn4MqHaBrz4zHuWGWcZWTAAInYrNoGMb9tjl+oqDdcSZom/g+0w+xo
cqnc73eo2FWukHuvvVZNgpqbFtQP5KvBXSQiMzRBFXQB5gau5WSDi7/+vVXun8Cm4LTHpOFE1jF1
kzP2xFDWTBz/JKWk0kB5VhZnetyL3aleVADvj9aD/61+pJjU84ZwM250rKvCBcW4W8u5mU4b3GLO
pkUkHwF9GkeNI18MHjWcQMf32eCYUBv7cGt7OIBFzTgIAENCCeFbBIwwMQx+202vIFYsG5z/W5Et
nOsShyxMnPI6KR7pfOrCIJdusGwGCHfbDxPWVkQr3O6bvC7Xv+sHUzHFQDFcXn2bcAQFSMvjfkVC
MC8wfTWltn/zP/NuI35DbLbNHZe68kaOyjCXV40xCoxUJNplNQvQZDoi1wddbpvlQTCtimkB04fm
KQN1tlR7wcUJ23/7oGE5r5ADRY2lCaW1BAKd12EcOFJZaqCq1GqLtc3hp0b7eX6QuJSE4hhbTC63
t/cwnw3Awt4NhoUtgL2vgKxmpWe5ier2hS90+ISIPhiH1mmQsHb/Rt0MM4XBU+GZwBo+EdHm2I4t
qOkvFIHg3tVz5Q78nrx1/BPgdPjMNnHI22bxCvTxM5KyzOd+wNWD9E0Wg2ekpeglSw74B1mcUXUi
tPNLYJaec4UfYQcH8lJYEw78tSAayCz6te6V9L0DiHeC5rUI8pPpMUccwt3QUowiouowHNJcj9bw
aHpw+cEsrIb0CsTXDrdQj/t6Jmsg6tmTO+gQpn0fuaB7rzSsZ9F1xzAAeJbtcFdwIbhVyg9PQdhy
mcHyAce35gvt/1Ht79m5zlM7ruCfHaL4reeFKI+EFWhz3+BJ8w92V3ITETzfYZ9+DPEFLZ+HW41L
J+DDS8iR+1DsefrJhlwcQbP42l6RFrYt6aT98R/3B7Fnpd5PbQ6ja5aswGF19jDVMKxrUbu/mUUt
VeyE6x8KUnpbA5SCGea4Y34G196tPgg/ZMaxrutRQWaUmFITDQMR4pbPIFxofgW6JgQvol0W6iNg
21YAT21c5cA5QAwHGhM1b/XqQKgW0y15iwlCiOcbTvdLUXV9DtT8SVY46T+0bEqsDETrx9D2KmNX
8f7/R+J5QUCO0uFN6CegecQ9NCFd+imzSWYqDwGdjsHM2vEvPNbxelboP2ad6gvNNTC6jOsnFE8J
Uw1kshiaaF44Y4NWVdAed9ExA1FmAr8zKn7A22rhha8n0q3DXBqFyJk8qhlyFczRzcwlxX956xb7
o/QRbiuCMdKrTEBkkkbqz9hdprgo7x/utCd6hw9LZ8a0kR05knLE8YBQ+pR/biI6Kf+/wT/Zhmik
YlAPQE9iwZn6vn4p1VuDiB0M4xys6i9frPsW9CYZN0824LY4IiYpk+bqXG9nlE7S9DyTZqKQVYr1
K1In+L2YCD/IhJPGbfIXCf8xeju8q4aMrROxpxxLcDT0eyEf3vF1B00OzeW4cHu1rj7scPW95Cvp
jlA04zPijKMkiTgBLq1V7mnfVpQmRsHTkyFdcgILHaO7GfoYtNk8sH3orje5lCujbnRtO151oyly
C5sFSnJwHGGuvL8M6VUBHLT1aeEzMAN1PYB2KEP4OCye9gvyK2DuSK6gnJV3v7EsKvpGyBkukrOC
nsbvUwndVV1FKTGcXF7pblYmLbLYQbz14Deauo3AwOhcIK2rAuaNsfTP3pWk1EdtLZFIRPYxXfju
dm4DbP1bTjBlKAItnAEXpFK2sIIeCeDTQV1fPSb23hq0I8a8wxqCMmMHDSUExB8/CNknyr+2sWlF
VxWiyR0vMbqsOWMMjyY0JHLt7E8FG26DymjTd7NjV9AaBM3qMhbIN5nDKVON9knRZc6iaKVYTnzz
oAYGOyLtGddngJN5mCxLmGN0kCjGu3eONOamywBRl86idy6DubpyakazDMuxC5SqF+Ct+g9aJlep
30ZODiv6Oca8DhjiX2RxRyBmvMh72cBNDMPSOX+OSbd1+3s+NSh9H1ndbS48TWwdlz0B0S4PkwN5
94W8mkxmyZvdtipPSK8mFuTYc9oJlAs2w/A4j7+A9hW1CL6d3rmb8jte0akYCTbf2Hd/AUEsxN1U
mSN9J5kQXwv47hOysHyF0oeMmsX+HYm7wAjCD/Nh47fFP81dIUVPg0/z/4TgD3qTC072ob6Z2Uc5
XvnBHigDT/FvI1yXWqXRMNw1oDLNUcmpIrKJvyzlckScI8x2igC7wDtYxBYcYE0hPwrIRrykyUk8
g6gg6EfdFa55LnhrGLMTkDtiHehL+DRxWMO9FZjRX/ZraDdveqLmV07CyS8qItFLxfn9Txrl/enY
Lm8UDQ9R9+XiOJdo/B0IjNa/9HbhE8rKJJToHpUoh55kUrtS/OAZyNqX1Hb5Hs9yb6l9u7dGYf2K
atyM8gCGwDpQFvpOI/g6Uc18ADPr+qYuUW6CTnn+x3i/pLq5PrKLceMjpOdI/6LG3psQ4O6L9UZs
CVRCt0RlexVB8t7IAblx140C8WEWoam+ClEGy+3uP/XJMPqXEnVa2MoQrRtCxRHOyarqw+ZjywDg
n7aYbyWCcfGC5+PDEokIx7bIZkGlArSbZ5tWwry6zLBQHVL9NQbKMm45MYfWhsPqgjC3j7z5DUhB
gHiGRxcIXANdLiIKYBxVEF0xufhYdlAOxnj/yjLXXTAHZpwoCZPYb4sud3EHgEVqCCY6EpH/N6+w
zpLxDQ23KUiMDK8XxZ9UddMt4f73z1iStCjQBgA44FPfU9edhw9qhbDMhDuGeDQytChqMBn9kxmc
U/CjDW4zOQkbgTA2KaubyJn8dSMmuImYrIclojtLFyUL6FfzTHni1lfhp0P8ZSOjWrlR75Y3e0ia
pBM5cUhdDNExKWKqTYGu/GLIgftT/i79iUxpCSDsaGsSGAeC4OYKhkOkhzglQupXzwynFkDMbNzE
Sypebvxu4shndGqfHGQ8c4javO2gDNs9BGcVDB8eTIXfrWVWiAQz8zXI9pGhBAPOmoYyjV8lx52x
vBDmUjfyaNbXphvOtQCVaXbRt1jv5EEzD3BKs2FHpwtpRWlzZ0EdLNcYyNPhiQ2iCDyTprLsatSY
ywOYLw/h9dA/qszOJxF6fNxi9Mqi8/P15mX0sAKgEl/YLgNAS7mQBotb4c/IYv+NIifOVf0nTBNe
WVGdfThBWw6QKd6SSi3h85QajVjeVlE3tleO1zdoVvKDLtAzQd/xtSkrsoYDo5NTfy8BcSldvh9x
ShEmga8UeBWahpYgSh4giLxJkFhSyx6iTLMAdieRHFYcDmLRXorLCQ0wImNIWpYcd3gnr0eDMnGU
r4WiacGF+nQwjIbAOHfNRIMFe0ELqSWcKw0c2QDpi+XYPvWI3IPDStThUX/nY0k9O3pWP65gtz+s
Cj2CKShkFN4hn/bhakFY+XJO89dmTB8m/YABIhjuAnUlRAs2msCJi2bF/Xp9kXk+YMPWSJoTaDro
3AJw2A/VwQU/wIA743zXrvUBUY+zWCxQNjM4mWV/GVpCOj8W0jP7sdiKwGxbhQuwjEgVFfw0YR4q
A4U2Wopg1Tc0rIGFYJULcdWw09fGQazJrX1yn3NdH8+2gWewUlmno2xk/luUljpiGxhvE1W16+Xh
grHn5f7ZWhCHg938Li2a0FY5ccpGhreX5kf2KMPS4amh6yfo25DEK9+PPnMJUuopANvMVZWsYPvR
HS177NylClDupJC+pOLy3uOALGBaPYWwXtCLC4vTWCS5nrniB0UnTRJb3jgpGWekHeFYKN/1fBsz
ILL38VPgwSgGAXdgfyGvXjxP0TD4VeZpIKHTN/4l7Z8e7gMuKdtaAa8V+MdFImNIC/eJed9LN21T
48nFTUmI7SuO5zGX67gJ+aYMCBME7bJA5BRYxStqjvVPNMEkhNGxNzVPcRwyTH9R0h9zKJaIiaxO
CgYdc0JejXgk2lGBodsfxj9HeSugOaPFlIA6cdyDwzgerdmMykLhYlkashqncirutCT8Nis9PW1T
qXKa/DgBVf7pXWdiLjXQM8M1w2nsfsFBrzXRx4BzEEj9NzyTwHxzamo4+pcdD4AqvPxEX9f3g9gD
aKgbBMrEN+5Xf/0ShIj1IeGqaH90c8clxdA5MwAvRnRhoX7+C6p1cy+IqMCVosfmr1hnTvBGCfZn
/HbBjLhAkaCdxZzOFxrVBKI9FPCxuP/nO2113TFgcd9DvOjMAqemlKjFLn8KeSEy+QVCr0gMvKil
NcA6Smj3WuRBvt33w1uyqNHYgPytD/lnlVwk4rCgx95a5CQ9yGIJ2glrB6L8POd9fl/nxUm/HTyO
lGlo9G2aWEmHoYlU1VuK9k/3xDDQZQgrDcXu9c7lqEoEzcwSJpOcvkwN0jRn+KkUvqfahwnRTASX
cCF1NEUcCfQtkbR1ifUTqXSJ0KQE5/gVusxGxuoarx8jKCrmY31RnlICaCs0EE0WDon57Keeige5
3AujqperZi9pl5cHSnDz6aJMBrVS27fWsqpcH4LKlo8rICLbQ9rwVZYBu7yegJq2K6gMcRlDh/tb
IhLp9JjDsfn5+EuGaHlTUGtjUu0esJXQTmiglU1C8F0oRma6GXcALgd1T052jva8JCJUpgW1fjbn
ojt5cOJgukhBHyqZPM8+P9bMVoky6zt45dHIO3BElTfXm6nRCa5zPAfAp339meZXOT9OkHFcRyEr
EZGiDxMgRBWhxXTrMjbCw24xHEZirxUKcXzJHOoAjP6TWNTklS8COBeY0LfRfaTc+bFItwRWj/L9
X+pyaneNIwewO1eWmRXJsH6IlpWjWevxyprzUaC5nv5Br3JLGIR7LOhP/GMlePGdnopyxAAjtqoL
zj5I3NFoan7x17GPfVYWPWGfWOy8zfNgo3AJ805WKus3qDqNttYEYYpmvopUXe1v7VUFu1gdf0RI
wR5jCLXiDGG+TjON91OFd0DX/OEN6yFeEfNuMU+ETduGgPmKVpQu02g8A2WzqXKu+0P1XQkowB2Q
xp7/q9aKJA4GFewwzCFP3TgL4K+dSFE4mWim3P+qaNiXmoJsbDwD7xjXJeVt6aipTnzRDm6nMnDW
DaKf+Br9b/tEs9OvcIiBNXHkWDmS0EcGbGozX9Vt/bhAT5v+2IJzie6U+6pq8NkzA1fe+YIv+Vpr
o9wGDswxYFz4q4TVNrzN1Haai00vlX5msMJIwnkFBoLgEnMQYyyOZovGTPAyGF6HtD5qo6Uck5xn
z0tJxyt7rt0diM1HsPTnxX4UP7iN0NvWF4Tahba6taAElSb3YDUza75mCEjhw7owiDpSttqWOdgz
GUbYHo9yam0H5bSjryNwN6jL2egkJJOuguen18hK99agwiwQODR+yI3dqXqMRkUr2Uf1kvM7fDzV
6xtHSVRj54C5doxlyM8rJteHZlvNsl9W4SRbLDjkjVQA3WIgew8/BjEVNpRglLjzs2pVF4jmYjbR
oA1B4jE0tql0SifOGEGd/X/ZIqnVb4ZOJysfKD8i6rWKAaqKNsrLGaJTvu4646a6MUiO8LefXVnb
jbuFes+EhxYEGxEZIcac2IiRORUnSnX7S2rXZTQ1V4JobplbWk49WtGiv5LaiW6nL8UnuNDsL5iL
7TPqz8jYYhj3ka/nh9MHV9s8pZ93PxGrwTAkUkej4Z5z9dJUvMSycw4cm/U4+LUlfL0pvVGSA3h7
CETD9Ix7VmSp4CkRqFl49xawflhsWRztgrtUgpRiKxP2/iNVjOSHSnMKRAf2OhnEQHWY+MNEEE/a
vQhKu13mHxSLX8Xu/6ElmAb6Tdc2Uh9Xp3CQXJzF1nIO2/7fiUnZlEt8Dvkpfhd+pjWWbxqeceQO
Zv6UN+ILczeJSwHmX1TWCLHtyhkW/+84NxFIej6wGY4VQnL5l8l3tRMqQ0zG7QS/bfHzbrmEV98j
4D39JbvqpbOYt0t7XmVee18Dx5w0ZJpPTDTKnWfZe4e1BKE9YBAi8s+70VzAziIEom82ddJtuK+w
VEMyYxlqFZxEklp3IGTNESV3kbUgoFRg5gL1hzsAUeasqWxP2HOfGd2UpkNg8mMn3/edhdvF8mXx
dCu2VRstSQ8O0x8pw8xwdRgtTACLRjJnymiymclROd4QLVQERjSMIO+i7jwUera1SRWGKd/VBpxJ
iiRS9feOTdHFDmXnbQMmW9T3UCMg134LWBtm9NYQD+3B0PhXAz7lXFZBHpEvpZwZe9IPXUDuBQf7
Ss+XuBJTvbvMsRjVeQQVqqEf7UBilTQYjrb+VwoaBuC6ZiWBsDcX1q165I92NP5pWfsLX4AlrpW7
reoxzpSh+Ue1kTN1BEIVVjy6iDV4CPOJWnJ1fzq6LN/3oLE7oHtxRwgqwYg++FvqMoYGwFRqFinM
CoQzY8a+Bgan8YcbbMQ9PbPNSkdYEUS4OMdzlIi7YMbR9bgmLvuls/JTSAHG+I7/GqV/rGpx99DP
tnqPPKLK7gV+xVrPNqu2FcJqerR1/YzmKW9SZNACXqAQTVJninTWt2ErX3O5Ab92RR3frc0qhlil
qLKf6HDaZK8pHoi4EqiHrtls/uZlLmdort5DbJDBsgKGs3/7dqcRBpVpyIgml4n6CnfzNBA1fsXW
7HmDoc4GpeUVRlNGYxHZ1acz4OD2x3Kdk3C/GminYxHCXyN3aeQnuA9pTvZsRmNSQo3Vh/fxmo3u
SW5o6WQnieLTEr6Ixzpb1yiHevwCgRVggtKoPSLtqxczKlu0zd2gYHl2FFRcxrpoxbqZ85IrB+J2
Y7/uOYl7BEUnL0TT9UJHWtwY7A8MR583Uo8IdZI8cWIUy+arf5b6Mkmpq2eE1pXavCF3m34uUmnY
AK4Rq94qr6acxBYRg2+dlQOzxjp9u2VKCpVDR/J3fFPpyljkOkP8Pz6pugpbEDMo9JuG6KdHgTPc
4KlzqNWBUP0v21XQ1DHtoRmgWRPWWk++2fDSvQMTD+699hVlwwJeMfPbRiO2r1J3jJ5d1SCgcpKE
Td05ZKP4bY45ovxbgrfQxgrVVKFHtpO5GCmL94jEFm3iaOD5UI7KdrGcscfJwW0vl+WMq+YqMKgq
Fre4YhIF/D3K4HZEGFEnC6K3rzKjBzS/p52Hp8fxe25bLDjqI5NN3cSn4v8+y0LHZYAz3G7PSPJZ
BEd4h6AQ4CkDRHJRPAkDF079A4YatNPryvsFNGVGW2odMwpWACYmAogWiyWc7dz1WbZMnIq8HoYR
VwD6f6J8DyBdbv1ndoDMphMMHJxSTcYWqZmvB49zHxmX6mqLdfJGyeIKvm8BXA+P09s8KmDrxAD9
caLLR49hyeLKUQ4N3hb+8RNGoWu3VN3gdlLvJFIqq/fybKX2+s6scxKcGM1GAG9UOiuFBc2DTpsY
nhhDiWwaimG1zs/a3mGkbVHDsRr29fGY1k8yosx2o9Eb+m8mjfbcW8PGZKjxWEW1/mN0WS2OLrIg
Lilby+2nD9jpfEjjir98pZ3tnVnpLrtq/g5bfaeyMf0rdf+6SNSNgZiWpzNVf5Pzb0OExqK0hx7P
gf5eLR4BfS8vXXndI7FlLj+mgdKHVDBVVIHq53a9943Xh1KytmjQc6kdhUuG8nO4GSprxzsAb/zQ
8dmzfUXF8WZ0SHs17+tCJhgDaKFCCq5wIg8YV3GQekTkfqf0znRivqJSbD/bT/v6oVPYnpv0zjat
yb9u1wrMbynOsBAFizlWUqtAfXuT9GhaY/iwQ8UU9OGEKvEdsoFLFZID+I24frKT5u+lZVN8XLtv
FPig7+LfUl89NGlw3jNRFrNGhrxhfNQ0FhbtW2Up/iZSPN9aQXxbgvcc1c9kKh30+DvbUNTj/+Wd
uRsf/b5tXeckEjOlx2vvF/zq7lGettEoIPuZ5NcY9e/se+kNvlA5jTMULwptykgO3qU1O++gRiBK
KwvHVNorM9vKT+Sb3CS4EWygub0r27tY3st+kdgSNiTlg0A6d8bUPO4HEmapg+LbLD741xwUOgSJ
dxUpez6tbohHn39DoG44uBu9qGAVmEYpSZU0AWGsCorHa2fXtfbeASDNI936G0DnXNrJJkxcFsy6
hVUlcxjnkL1sUveVCSR6dZye3GRRSYs/A7DCVTP+KaNSOTc2C3v9WT7XnDA7A4ZMJjNDlfEwL8KI
r35jc40FtlCazM6hHdiJCKaxLvyhn+gurf0DmFfFavL/cYkfQkYXiPWN/XbGSRqU7NXSs1eaOuh+
xPNqCdske+un1LCj6OsoD3rWarj6CrK25okHh4O9linMUerFuC9pyWoKkWUc8QVJ+UG0nOhNhyib
6o/6b/iy2tcMaiGhzxDqF8BguyX7D2SmWawKSUucpFRl25e7z4KFML47qSkOSNCy9HOiM+Cmvdp+
pueYe/akYsBqJhKLXFJhcI8kS3FeZ1eGmYCxPUx8zL+NJEQ530+HGpRhIlyxCCaxwxQKLdaKD5yq
iUa82i245CeKKdoKWXi6g+9j1derq9E9R6BjHo0Mk89zRYpofymlzkbUmFWrhcTjbpduoZJ5Z53W
nZz9qULvvvZTum+HUt3OoRIDzdxKkbAdFEjXPe4i8VXK20ilFNQ/bWf4JHa2nlFmmwzFgKs2LHWY
ROVQzlcXHLkdPfDxHa6R6zrxErz7uIUo08yTRtYJkDG66jlSsN0YXH48IQnYM5KAj6NYBtv1/Srv
cuVTJfo8bRUiNGcHIAFtK336x5PrtdibE+hy2xRt+NwX5KZJEfpR5IB2Q5JnJfrHLRNYeNenoK6J
wyIC1n/s7T5q8xiZ7wyVCgGsVq9V/9WVRrAERVF0xDTqRHEyTTk2XqpMLt3yhRYwHdmlYXqQTjy4
ApEBFornjlAKVBugIpLdc7bHA8v8IaqrpQSO/n9ETybefJP3MoKUIEfm/xvgRLs4p3LBlw1YGHYl
akZtMsL/iQ+epeE2ouEsgzwoti78xdphvf7ZVQgIpeSiOV0GT/JyTb8xoCuzSqyKDJxujggH3N+G
YPJaTP1x1G6xKTXBfZH+znGpz8WvdxoCQLJnX7BvkYYD9X6EFTHj1XZ7OULR7fft4dk5K0K3IhF0
YED7ztyFquxHQEHlX/QC/83DorFX99KORJqcocEIbft0c+u5GNI4thShBK5DUwQhhPzQfvXO8AbF
ZH1VDYOBTvgYdCxf/XocLwWoQXanBLyiPYDNR5gccsvzGjBYxt1bdAAT8zWkXkHxAGsAz9Wh/KNP
je6UQERjUsULjFO/xYzFJMvFZ7U3NgkbP51tKB3UadYLq8Ddv8OsXaEhbCeUIdhQ3toODy+RaBXS
NCq8WKqF10HCAzL/n6+IJyMxfDV+x3A8OSzpa2TNg0SrXyGzhD+Rhp7pSjH9cz88tegxDT8vpPEF
Sdu20C3Ti8dzIxQ7PHjL0sD2Cf/KdzotAaieM7wSU4DLjOp8/XQbbesmxTW2EIVWnwe2CAg1kRUL
ecSR7S89vQdslgw8PjQ0ZxxI5V9wwM0EoUPqZWY0Gdobdf2m0roWNMlGNd+J4azdVhKjJqvkic1v
FQkj3Oee57JNWRUwVLV7PGCYuhjqZ+srrJKE4DEHIQrlVUHnoodT+5+bsP3VjkwvJVvqARaPHycY
r7AYAsXS73JLhNeuzhcKgMDWrlUo94l3/CZ/pJiugeuMpouyze2NDnBMNtTugEG7J+jdTnIcs60R
cgpaJfjJsib1NwIw+PbIuVGqSRSjDu4m+NunbIDc9N5+f5nflmitaMixus31eBjmOgR1JycLowGv
SGPDm+KVuV3elzgfzXKIzZycdp0DwMMZCjq669D8ov8cimv3W8gVvu9AYd0yTJoaIcVkrYMGZCDH
cbWe3u4sSGOQIKrAdlx0Kk0+7ujQcNSXN5r7ujono3T819r6WoSk3RK0rJTjDYjsH182UWN6DRmy
H3JHorg41Rf6XhBklA+hjd3p6QLvkV5Qb7Y2qlDNtWx4oyXxRGprlZusByg0xR3beWNZ/yYnSvZv
6PELb/mbQtPVfv/8NxfyT0kF3WEzko2RttTIscPbdV48rjDpxXWQSn+dN1+PwQdiZIGWrsTujBgB
MfFe0YobgMld/Ag+CQMzczMDTP5kICXq15dVubWJqKYa+0p51pDFaN2UJ/rGFnOCEEVY7dPYGR+2
v9JbheZYBI+g504Srul3n8DTlRY1jwIQBGV00QsgrGM5tWVqwzdm+gbT6VlkL0TKXQ6BkYudhJGS
nhjxv3tn0Ylk2lthTTRugrHohDQDrkOT8SCWI4GIZwlSAw8X5H3UlX7ydohwFSokAziBIN/AXGfr
n+csthWjIQYjRA/L6duqtIxvTrY4iNyf78+v7SFk4X/0F2NcA4+zDU2s0hMS3MT2AzXt3SXSi8ni
xyrGzqDjoRcA4StfQDX5wkZ+XAv+sTEF5FYhtyZ07yYULVUcPcTIxY9ZrrIpHNoiMisk8WgWLkI5
sJbj1BXONJXTayy57M5qOS0rnAFrZIp0mlxL7SFiU4xrwMXmFuZcxkyyBRBHok7R/8zRBGEl3Je0
wq0Uxs3Wb4k3HDJzPSBEaokMaHd1T4hFbCsh/WsG63hV4pqAvYNg2neWKgw+cE2IRdUEWsSiqnjf
RvybvT2hJ08UbM5xysmsdtTssR5/V3wrYV7lrPheJVY9E+znYIefNpmS6xB1XxJ0YFz5sjWAW0Xw
aWd3vkLmxo+aBh1P0HIrdGQ+RbhudR5VGrQfTt46E8OQ5LZl1UIHqm+ZlG3B4BxFsm8mnTmouuYE
yz8+9gr9yZzD8grTbNVTuZKrJxIHkyjurucVkdjUA5JxPF1rIaseaX4vhXNPxRHtiHlLTkMb4zYp
d8/Tv055z1slQQerBxIc0dsqGnanKF+xeKzdx05EXXnDxfzzXHKkjPNCAlg5N4QQp1hmSlfBGm36
PciAGqSCAjyiCpOAJCt2pZGH1PuRu/ub96FMYFedVL7CDxF9gi4SeVR0YryX26KDvM3Gw/PzTRxR
cPgOllgJWQ9tVReM4/Mma9FW0hQ6jMwQYaUL8hczr0xk9NvfbZIcO8v4KuukdDx0qXbacoSbGLjE
t6Kd+uZa90f+sMYiukl8IUOQtHuIZCvP7gO4o9VXjBji9ylKcroM+ZtNQprj42Pt9c6hBQjNCWeq
QELXd5+656CH/gbUM6JFl+NL3yJkkTfzbt4fKA+ShQSWezcBze3LKPlx8b7ohvHFuamUsqapBFmK
Ws5TBpTh75Q4rDxmpn+DvelNXM5k1wsKR0z3CipOTKVEzWq2twrxVl7lL6QwDym+wsIPIzDsITSN
lF8ubLw7PGOYScVoy3uH+8u4K0Mdv2qtB/2Z57rr0ZaWx5+xE2mi1OQXgv7EmmUoSU9O+NCAnCAg
ryDgU4oIQ4kQ8eBdF71Z0uB2sfrwn+rKOAjfW2tu4hm7Gut0NFQrp7asqJEqpV9wwMGVTsKoWrUH
KuLT4ko2iQPPv+puVqORMMB5kW2/qnhUD2hp/W2qjRBZ/4z6JfeZrgK/0yYwpRcP23y70OPiKyaf
i3bkMNJaJBAOeKRygyoJMI3WUB0qE0M58THo5f2HEXKI83hKVT8n+ifuFqQEccv1sf9F72GbXBPN
yARZrdfqhBjmp58pPNl2x8LWIbG3GCzoYx9/Z/dTWNuxfQMoKbhQPii3LAkU9NriPlVEaGu1PC1a
/cy8fQC3EU034xcyxwErdEjvfgyFRBGYfTU4smewtHPpRcuJDaLbOY6plYp5JxBU3CBjjaXIZH8T
cSkXmMfGbfK/bZYC8NTm2e45dcebompVVBGv5X4xRedvWYV0g4eanxFkHq5A1nh3e87tT5CS4X5A
CHVtRi9Edw6QTa2laiF79bc6bI3+OUpU67C1Ebza3sf2TihaDIycStkM62DdfyPesdmEe1M/2kKB
UNn3dnYzUeuAoXK5pHPLAcVnWWuRAlasQGTDDV2wCFoMWdQV6flE0qvm2kAWsVPinXphFa8oBied
nkRy2yi6+E1FR11t8/w9S6msDUFVamPKMzyiqEyLzoh3goXgR5WAGwHELzWEqlLSAv4Q1JcYs8By
sWc8ESugCqcAgYg0yQCsPL/6B5uoNnxWyw2W53ALZFCLEkbH7npfktlOOLeK6u9EFtdiTME/OF+t
zkYV2jFk5ybz3ZbcYolrjouy2OK49RaG6jFq+mZP+nRgV5HrXuZnwCsoqHMnnMD+o1/kQ0mgIdq1
DmN8QfijKdRCCp2VAph1cwlq+5RtNp10ojQ6TlyMzj6OYUMg9FjaoMJCY/Jme0/fKGBVtsrxHwnB
NQnPfvb0nppHJ0WZchr9ay4hMn4eEx8aTfFCIliuM6XskKd06hEJz446a+4EqQkirlV4Cn+ZZUH3
VU79lxOGUfbk8fdoSbXqJIiupImGe2Y8zUPLQEeJair4IJgkvCLbPTK3PrG5Nc60GkV1Imr0ESxh
WouIr4z6xz58dt1RMEG7enk1msEC2n0P9KnAU8+v6SIRPkLXkHDXduV3IOm8k0P2bFbDjYUFL+yx
tsIlLBJIys99yMgUUfmxuvYOTttxyzJ2XHMpa6YTSQT6EJ84smV0MFJY7tMMHx2euzn5hLR9yxc/
vcQrDjQJDpHHxPbLXWna8EgHqZ/QRbz3yq/GEYy+XGesWnmXQqKfWarzEeQ2o4GAQbpXYtclWcle
IuOTKPgeYF73kmbOniwMABYTMIdA/KN5nc+paK+g4j6RmlaXozs/r3/aK/eEH3CxCjByafQaJNeO
EKWKHRv2KCBKBW53Q+iaoFZdYZ/zaasHWzGuB5Wz59OOBrXH6UNZ6FotKK0hO8yIhVjeD2dW4CIn
1E9ARHDV6HkCspzaogBlVaTXO0xeg40Zt44gzfU5+amTo3H3dVKPg8ceEmcH2Y1G6x0kClvBc03/
PvUXFiHr4ra8DtyLTvh7VRS2n0UenVWRfb4jko1opovYKVeTeSelbPWul4bgS8Aof1cdrn64SluL
Ss9A+ZgITl+2ro+TCx2vFW2NCq2MdPEVmYW8ruejTRL8jp+dggSDPyKN2IKRXL7P6wNLzXJNNltk
nUh+dtm0U50ygiIHn2H5HtLCIdKEg1Ni6sNelIRXHzDxbXOe5UNjMB/BaX9L7nkl54kbZlT58U/2
tj+lYqUJaCUMGC5Bv0wSxIhpq4D8e7AG7N/bWtkCnn+Z0XJ32iVQDc5t06KCmspiiqTaAtJOHfn8
n3OByM1Q/AUBcJJD9O+jRwNXfyVslm5A2es1soZ1WRQ1JBIDncsqPnH0uJjvWcwfo53Ykt1XfPlk
KlxG16W/mAL6qiAR5p+gKtB/GsX+jrQm88CCW6edAW8DMyxoBgJquPX9+9WJxQZj0gJAgPOUe4bp
j9EpJaTvZrUmPk3HL8eIDXm0UqMrJCwOZeuGFAkyTcV+b+QnfFQaWPIvI3ucSKcmGWm7fiFVph2z
o4OgOv7AiOvDgt5dgVZ5rPI5zwAxclA5GJXGfdf1gsGDIBzc5q8OXsXFqe38IelcDxcEWEXrB0Rm
uxbenbqnipqaZe2cCOLWrdcpqJLF7n0rY4/3M0tTWd3weglpsKj6xSmJXB9Q5Q27BjlOt2j+qj6Y
2mMiPQbvHpWFgUuFHyWb3pw9B0LKjzGXvhuGZVdoHJV4wXhA+x2BIpfdN/LDTfwHMvyp9oLHCxlj
h7q2PiCKCamGe3dycspbqE5a7UHec//xxRu0xYaDeWTI/1Yi07faEOkmURPZ0Y3ZV1ye7i/wIvjL
0h82oO+iz10Aw1u6yghSgVC2lRafdxJCijAF9SqYbuHksZ5smuP6cs0jryQqHIyIF7oKhHZnotYM
op29FHwe72zIE5v5Dwb6leaSfHgPvsMMF7JaKIeUg0KVgpUelwGQRJpYkQQHTtd6EdujB7Mh70Fe
QDw/bsWqHmGrEqVx4ii7k40elNeqgY/MTku6GNPEW83cXZruhru4SeUqUSGAofxmPern57P11ur+
cG5yYgHmr018fKOGznfnJJVLNx5BVVt2m9ZsJNlliEVPtC4trJucqnFOO47Pg+VN54MkS90jwM4a
lSX7kY9PofnrFhy2w3k/FdsIKTLEgezQneUaAj+YD5sSIdmcQMuG6CSLn7Tek0CNEpcGTWs6Opjv
gqgx3KSXuv4hA2uB+LIUrI/hoQq+hU5G7jSmt9JAEuuGqfN/U+WEEPbG2ctJu2MA7Wjer9T6m3a5
2LHX2uutMCymHBVaJ2Xt7MrpuMpCg3oMtS6dXnRKUghcDfpcwtPokNZJPvQMG/RARq4c947AqVcQ
ELGFF12cusP1KpXUQMu3VE8DtVpwjksFi3EFo32AVXqtJFHapBSPj+C8sbf8dMr2tcuPygG2TIP6
bFtzPOM4MRykUa08FsJdz2Npsw3TnEvlb88OLnv6lQmiwPGJTI1gD12PIC9k44Wfx95spM7NDExX
J5mkMMwq23EWKDy4KJULV3JwSfNYedpwt5cOZY6wTociEFh80gaJrMTwRqbVvwFF4YUUWb7wbQ05
vVoYM+2gPwO66iw0aiwJ6wJ0fqq+9nQrQKYgYec3F2ycvCn2Ce33Evx2J8CiN0KkwBZcv4XliZ98
ZCHj3cjG1V55PZl87fGLZBswoDkDi+NNduTv/2P61ycCY8kmG9sKjmEWqHJo+/RTdgkqs352kFmb
QkJFmZ/RMllSxG44a/3PysY22ObwOwqdFjbHYXOGWy87XtuG98NWrQmO/RHRQSkJGEmpZKkTD11V
mzlPeSEOJkJ/bzjRwynGEkp4mtASHwkal0zoYarLI0dwK1jAf8pPUgMRBsx+LXQaz9a8NH4Ow+RC
Y3f+002wAxXZnj2BlbfNi4i7Wke3PR7pv7OnOzHm7b7t8idU+xTtVqjdNwNlTYX3QzR0shcElojM
IcBWXTZnHED/pax3XxNoenyW6baJIzl7k2OxucHoJB2Lw90O1eE4wF1+JimTVxcGwjPnS2vUxuPN
o/HS9kXtVnjxKU7lVyxMkpzgC+czgARWzB1vUn0oPSAz05v0PFYk6KrooHlE/EnM1UdBsysjS9UB
9QAdSLAhD8JU9ogjatAifkLG1pROn1gjWjAb50goOUM752UPz2MmT9wKRZYg9r75G0g9+9ZBcsUc
02gAc8RR8RWYr6wR1yi+W7zL8TDzW9HwsIoN/fi8A8yN6o5+9ublYZB3/NEE/IINCzU3ROjdXKtZ
yVm9GchvAuuri0DOyeTq/9B/VpWhAMg0PIx67zTATkI895v4+WE7JnuCwfPyGhXknhmnsofSjft3
HkrzQmJMUrgWfcU9lXOhYoyhfB0uSebFCS1tLzSPH5mz6iBscs5aGxtTaS167Hbaze5RFLefTDvo
W/SGyowmYd0VklBBrWre6gbpaJWjur7D3UqUqmf/RotWwy9p276UI5JuQ6HrqZFyZ7LNG2rU0m84
oUqjG2e+SMSQaINNbyucH1gOTqQZwO3PaE/5ABGUWwFM2qc50G/Mp8Z/Ob8FT443gHnuts+Y9O+O
6qA/BUBMZ0/1t58GQfTGa4esXkfsDXXF2lThtgG/7YvMpkkLy7q6/0zxZ3mtKpudGERrkqXdQJzS
H8a4xMWsf7mmnAT/pRTZJ+o7S134VKmkdjqvXe77RMD0ENCojtOwR6we0NhEgOxQnOAZ2XT2pCCV
ptaWAopeyrQ0kMOzJebV4T0a/1H5dCm2/tVM8PcAdhe2c3jx6F6k6awLnB+Hasm+nG41H2NYRVSL
8SPrXZQVKp0Pe0QMHhtgBQQ82vzLTLR0/ge4mK+uTl/lFbhLV6c7f+MFQQdaht1Op1XKORKkWL5y
ta28YnqRtH/groCEkRqfY2T0Q/bvJXXwQHqwpE+F202r/4ziOKbb+XSCgfaJuwiWMCXrDDjTpa60
uHBeKuGDoP+PTVAerQ7W85eOxYdpuLzgzMofaJejuwjuZ40yv21rHabGsO07Pv/kUYRvEhzXvZC8
BimKpUxxdplnF+av5a7DgX9r19FxyQbIf/a702cohcsvJI79pT3v3N5Jn61tAji3c8n/UUCS3Hsq
NTp/Q//1MGChBCE/jYi9nmVtoR7kE++1x5LqyyQ07S1qvjM6SLSzwVuI+lebj5pLuhbRGFOKknsq
8O9iq08cTqRc+bC3m5KurQzGfBsSz1bNGM24FHaj7Qf6fTR9Gz3JEZUp4vRRgHveorvkTggyeQ/f
AEbJpyisjtZmAVu37LRo5LpD5mzc5D+XT2jMCr1Dkte5ZzgAPe63AzrRuZTKGOG5T2QLG7aFenti
31u57BGxBeo/TpthPk4t7TT5BQY1PyPZ/tS85ZuCxm8dVKkcsUgY5/4zJ7/7AFWIXZNKmCL4ruH/
XyIaoHB61wBTUeoTOLWt4tG2sHgllOj8eQ5fOZbYjfQVmkNyIWUbAyExZVGIGr84peMUYU4z3PZy
M2NsGDsG0YsZqTakD4UAL4gx4g+4JnRMofIZaQrUVfDfbVo57wff+JYTAHFSluVE7dZF4vmTf/yp
v3wKQpn6pUckDmKxF4NlPu98ztDkS891r2glJ1CsRQd6QVLrg3x9RIOzY2hWNaZMwg9SjxsrDia9
2/2/8BXs+ubDZIroDwA5hGnyIuV7D7AA5JBJE6G8Aif8R64nA8aXNmv4Z3C1G6MDW4RfGrG5Kd3Y
wgW3/Xo2JUomkfkrnIJ0H3I+X6f8AbpBi5uHV3MewAPmJoWoJB+ERdajLk/7cn0wLh2ZPNy/0082
AS9fOX+ROWA1MKuV9FaT5jk5ba1YMmT8Z1hC7ShfacOGZHaT7w7TIkuSWuDKN2IMbP1AdXepg+w2
8wBwSFWo+rUABy7WVyFWhFuAaRMzvwr+TVmp42KaEXaPVVm8rCWSgc4HyNsmxQTnvZidoOHXw5q+
53Gq0AaMprGyzVHySpomr17KhXu7m12y6GUCsAoHsjlD4K0xSBC603AGlPkBl80tlYlgw7Xd8u1w
lNF7nszLbh49lFYsLWFpZZLvsm7fHLOV2cVIukTx16YilomlkEKbP8GmeHHeMHQCy1zV85jO/9iz
U/3ozeXzsqsy/G5E5SYNUe3Rd0luyWS94dvWVbLAgVqXzjPBf7BJO2ghc3gd9l0HdYg7OAjzXdNT
nnd2UdVLqCeMf+U63EXj87X/OC9cdVN0jE0AxCrbXq2gMhhTTq9aoN59EOOKDZ/S79JhNF/N/L1X
ts6Tav8pP5o0WfHvbk3hmudnbFLcbONmjh5J7df1selMS3w8KEdISvmY3ZoIJJ7w1XwnWnxS36Zu
actlhgvIDb5rIf6H+t8EZ+uqX1tQSAh4+aFsmIwxpDz37e72ag/E4d/SCfg+pazXrQpj9pAkeI7H
1sJhZsZV7hiTGCelLgdHwQsbJPT5AYEJbr+xBO1bHkmgD/1qMVZeNoCk/C4kcqAYrx3utYr9MWON
hBnPbfLvWdjfPb3WrVcEpGj64iWzRLJcjqjutWd9UkrH0wSKrEC3lK9FBf905oLuhfOLDsvOTM97
ZT0YEcoi2f4XQznEQANVxxlBb91kyoH7cNH4WsxtbItPDm1KgfvWfk9fDriBr1q/LxIGOTQfVwGh
vJm5SYrsNRJ+KGLsQ0OULs5D0J3LHNe0avinLaSYtDERCF8q3yvCFWPAM9+Wvyi413oHxYzJjnl1
+MsZLsdCZTaaC7giJ8QDJV/Xv7xAMM+r3DKCiVJ/nRUmfXBIM2fz18/aeMA81HETQOe5bKpQzF7w
j+ObNFsIcI7DU3I7j3+O9d7gX2exLUZfUxwAcGvJgTY7/NJRCTUOMtG8WFsba3n3jJ3QbG9UAmSd
DvT8xwKMDrTqrvLAO+foIO7H8jejIcysUEJAepY4LPffxyUoFieDKt1gfr9xN0fKA//uDGZSUSMh
pjAmGXPR/OLkjVBwgd7ye1v+cL9RytdXquylgj3IxzdyrHFrNCVyNXqaesWY/745uEjrB7ofW7B/
pz5Z6sPfvjPfjiFhIJGRBIZwQfpPRTcYvyj3GABh+WVd+hhrHx1wcuZRGgurOH8QBF9yXNcbF66g
i14dJIb1VZi930Z1v9MbtTfglgwDgpq/6mqkeqPRzCJAg/9HKBAb6vS80qQtDHd53if3wiQAoom8
OOKQN/C5V0Fdxk2R6Xg6dmOflfEx0sj5X0X2Kl2r+4sjy100FN3epuKfjVfVY+WxGAt0tgTc3z/Y
ZeL4k/Z0WJCx7XRCVo61w0m1h8S/I7uCM7u+Tu/TBtDMK8N1GwMm0ItOfWZwJXZOMfVf4LWrSXzQ
x6hjVakHMXg/XsnfUAf0htPGjse2ceBi5rQO1TIaMiz4vtsYtj/z8sZy/c03BF0dk/dRqFNwTyV1
AWCEyNkhVcsLwF9GEsY4YnONzYYczmyCn9w7NEMwu0JlRU8HOhU7qKQoMDUXhycDvvIKSpw+PxWO
d9IY8fcrU3QJ1mxj2I+NgTgicG+rANNai8f35g94R+xzhOhBVF2VyE2JxGqYA4CSBNFwZXPtTIxf
UabsPyXWgjJYKzva1WFmiVpPbmjBr3EfFR6IcXoNPa4nR8iW9G9221n57mOgQn2n4Ajg4IXSG3V/
nbaO9IWSv2ChSvGDm0S9+7i5aV//6ZYtaruJWgYvcYKV1PnNdy2WMFHtt24cRpCEAkaWUFpi8RW4
4QEwyDwt6IFbn9NPo7QYUewpYAudY+gVFpKAyDqaIlbgEg+QUbfeM4xFMfQEeAY0NbJ07p9G+a+K
eFgyktqE9/qDPWLBwkI7YjDriKXMBvxD5X4Ky5G1qYrA7eCAg/x0lwkQZGdDhXBF6kUtqHkwQHmq
zZmHy6ZNwIH8D90MW2Eyr8H3wL/ULsZz1v63aBQIYYAuVT1YhBK2DTBPTzmGpzrp8MHM2gpMv4AH
gWGwssfsKoDuNXXjDOWCzdLYT+HUYB4erp0tRiP6nMAawloWGglkMwya2g36RXfM5vqwxXkhhjW4
5rEypJLMQTmrLeSwaYWbWqvSLUO8E4JNQsoMdxlUHa2uVCGVJMEJhHZmztZUF3VvU6gjMlJcHFpL
cp5X0FxMFa1O7+BT0n3WOfhldhiOVhdeGvJSsJaSkHFVSlzzLmK4+2j6qLDUhIgmc56X1vMSum4F
twPgvQg1riBwbAwSFpFZ20QttS+4rEWA/U5HEQQZoC/NKgcYNjDFoznedJZt7hF324P+04E4WuG/
RD03m94deMoMezGsHcIKaH7I2OA9Yvrgdgfo5fkX0dj/+ocDtBS2XMwqBjqEOLAvumJ0q2CGTqiT
vAsAm/D2Su1/Zljd2EnVu5DlCxnPtRL94QvncChM7zC23krA76pKsFnREK1Is8xyqZwBErr08Ytz
61QF4vNmX2QXvhrbAl2osZeUAHGBkzaOv0LuY/j/JE0ioM31krkLHd96NzxLdfAOlS3BZ/gJ/eYg
DqPlXDsyP76t3Dcwd91mQ7PwnmoepzXvy0vEcPaXkajaAJ6j7bHncGm4lkwHuA90vZxxwNXleX4x
6oL7zOC/qvpD9t9Gb/ZnOHC0hcPadldGcm/JzPwLISSssxXWtp3jU8X4ectG3FQnE/CbknmfjUpV
/IEkF5HFaVAgOmxFMtZ/6ri3ixfpHETcag9aW2F72lkz51bcCdspviuCZez2bFXpTaAA3weFkTs9
ZMaTE7OOXyFRmvVcDEfQSKNUST2xbK6viGNpwGIr2+ovfRqwUMuQTCT1Vh/Yxq4a+7ULtgF1JNXu
ofLWahJvngWi+PIptApf0kJBmoYWNmFWQiDef3oL1n8SbM0hV3+f72xcA3iQPywf+IUwA+TsRuvh
witCitc1LTJE2MKyl9J6PLBmDMHo6EVSo1A64+JwqHjFG+W1Gsz8b+Yyp8u2JfvYUqTNOfZp+8gb
iA0o7udhp2HkoehjNjbBArBzE9rXUBhnD7tjgyIHmf8JyLfBqs/Nqg+bcwNgyJnx0v9d1o4NxSq8
+OZhrqTYgPw+lF9QmO5XAwb8snfiGy0Xx7mK6DVTjlU5y4J6WNSpw2WgPLokhlDGuRgGcgwB1WcJ
Dhrz2coL5kLaMv90pP2ZKklyjKV6HmZL8LPBYI+L6eUCrbxr28ejazHLkWRbOl/OIXO7KHtePOHT
v2KjA9FsuSiUoOVyhKXDVT76KCzDNgivfWru9tPKxKGdcJFzSJSgW/R5TtvcqeAxNROXHGt5HrxL
VHSwPQmygzFWCqAQCAdbuY+76t8934RUoxhxq8cWZPPTwd0w4AstfDJ4KWm1PEGuS+qio5aC6lFU
SB6ampgO/mNDDwVs7PloXea4XJl870seAU0oCck/FLLxoiQpYLwLIV6uUfD8DzkyXhldGH9kaUX6
JatL37ZPDo07tWR8rhJpkJvDtVmeq8D0EJY19pTeLggdg5V8NYmldE8Sv3aPaArmuAZTDqx1e+w9
FThIhhgT7+3qQCNVsY7Yr0xkfKkhUKcABXfIT6xECEwNoPV2UqZ0XiyvdTzwTJAuiG0i79C8GwJI
2bVqIYmxCMMPi7m04f2gozsV+dNN0tnGwaSOeHjazrKI3O9tOgDO54x54Wi5mTKbSmYAEwGqtqB6
CAWYGIRj1gP1y1mm83mQT5DpUyzcFC2GZnavi/LHRk1G2wfjw5yXZuKNG+UoScMsIdUXg43s6jvc
Kad0iGMo8qb8mPTnhhXuNNv47I6RsrFOjOmzc/on6hbtF5V5uSqDrCL6EQfSANso2VlOukWPqXtV
1y3RiSbbiuq1I13UYxRO66MuSDWisifM9sxlvzYe/hv7rVWlce+5J7NHB5ihIGoOLKK3QCVT1CyA
zgwKs6yGTqYUafy7tSS47SfLSZ5gs2yEaPUvyBRlSFdZeYKy0gcHZxIXI8/ZDXTGlr7b7qgXdUJ/
kJRpMmlHmvIpl1hyXPn+RTTYqaXNxUB38OpdME0EXBtchvoEP87TcRJHmbP7FiW6NCV/5RFya+5F
s3zPMHRy7472U5GSBzW0ZJdZ3xOXJuXGdCj8ggl/NCGzRKah3q8KiZiMKFyaz2qgM0fVYDVVnXaE
0VQopEQJetr10Vc+aadDoNKy4MWae9V3o+rjgDQCTqDrXEWxsF/teiZBk4nVKXESMNR60V1k0bSV
UEOif12RBhyJzFGoucRI/ws1Xoobl2b3HafT5y3pjmcGj146bDki94Na+d0YXhiviASOtoDDC/fI
ZpUFymBBmQ56ExMvMouO2I3eRNo8e2McR+hv7R30hhwjEJSDUTxIKoTaLxiPlYkkfehb79UGi68C
msv40f8HDQfopx5C0M+Zk22aZgR6EQ/ASugZgaUV+v+gLR3TtqIO3TpdOHYY34Dff/kExiHCocwS
L6FmM3GJftgPxHm5lAf4QKnJY7y8zwlPHI/k/0L487tJBdOQKHp44f+Q7OwUvStY+aB2zcPNEAQl
dc3Xdmq3gvt540Cp514xhmF3TFMI39npJt4OIgf8lQFpst3faEsbM9thQwxMJsrAbMxskdvwVBTi
w0ab6iOcNUS/u0XBVIzMPZc5Q4ht/GfXbKBNi3uGfgY+VM1D4QIo/JQujRsndOjykq0YZoaUZy/T
po5FbJosyMK1PFLROcqStlLXkcdoRGwg9elkTUVlIkesgq916YX6mURuSeZAC+6riTc2wre7c42F
BtXVUDt7CD8Prx+o6DqNFN/lCkFZW9v9qlNhL0EhGUStu8p1d1qZFJZNHyloq+4sh48zMSfdQbh3
kaEkjB7KGuYRsi4edGqzM77vm3Gedht067/o8tC/HMnjU0/6Zvv/3fhGLeJFEDo3SG1aJagiT4ql
oNDxzXuHZ7UZv25sKacRejRHjb1koMTUAuH0ZQ0OqgSTTQdtuV7Xxec5jqRDCVBrZwkNffJE3gkE
eA3Ct6UXK8ZJkHr3SL+soEytLUexxQVLUw8p5th6bfy3TIsBLLm6RHPsCsnjQqIzcJGJd98fIqJk
btQNZzDPwEqBmDE939F5NEJdPczpLsTgaVFUWNrRe6b/DlwwfOsjY+lqk/m285HdZN7bixK261mz
ApYPV63YZROJJlyRsDTl7U95407UIqnavDzckA5Rkw0O9PQ0FNgz4mZp8h0l8ThnjuBoW3NoYCj8
CVsuQYpOajCOYNjJEhuaSLEhyLOoHlpmli1GinH40vgE1tBs5gnfhpDqQDJ9QJVZR+CIWp/Ri4lL
PIFIjsdKkAm4IueUViFHEMuLH2frtfF6VL7ka5/v4g6ZSdDbIpJpPoIyuTgmL0MRdy8pUYNOmmq5
338fjOEwNDKqw5mdEga4WTgn2MNjTJrtL2wDysqree9KlRDlEd/MqeYd3FEMeN4QGfQhgEQjWNNK
GZ6dj62k7MnulKIhY6BivJaFVors+ZlJpTOV8h/1mJWriflhx3iWB0Nu+DbZImPGDFxRFgNg3k2A
BoXqxcyS9FEdq79tC6w1Y8zjb/W3YyFyrEyLYAK68qBOkn+We11UtKoZiPi5kfyVyUFjf13uQ0Pz
6nNnEE8/qL3J4UfRzJgugAHewTC/rmIegjR2ePtMvZ4ZKPqKyjKVWODrDRv4IZH3m9Xz0jsXOG4H
rCuRiuVBmb4W2mXsRPAJ2v5nkw8/qkLU3m06Avp9D18HOJVE9z1FTj877mupvr7yPBdoPZn1KMIO
qHKth/WoYQdH1IQxDXL7/CkUB7kVCv8F5V4apXhSkj/6IKaRQE6VfilfL/dTH1HLYgwSnkJU/Arz
mi89hci2YTPGc7rgb1Md5NBZXcgN9gRN/2oEzHknymwCecASBiUOuasqtZXrmFTnMRqs6Bh/n0dn
Fv7RDIalwm9jwXkDHkzf54UB62HN8CyazdBPlHxfYE9TVYKICd2lo1Iv2zuoFRnV5Na0mLNbM3Y5
ennZDgeMMtpMEd9kFeHCHljdQvMCJB/K/EpV7RVd6kyzJK2VT10kkz05l3p+ZZ4ua1Nm7WmkEJkq
Uc7j974KtmRUVtBRFXC+TsR7JvqdqWSQFklUu5/Do7NZY7xHxYX7DZJgUu6FRentAAa4vEVmH5se
kP+VJ6k4GDiTD3/19tiulYI+ICn0XblBfQ3QL46l2SPSLtm9YsK6Fahb1PevFv6eQX0skRQ0MzDa
I2+smfbZ8RRU4ZOqmjei7lEfLhqMhvdCtD36lZn8kOVrUk1mH+FdmJ06w4vfh6VeJmH14+YAASow
t6F3FhYhH/k62ym3JryVX+WIUMBSfgfw20clC3sPSYOjWbTWYLGo6R90D8m7mSxv2cZKgB+vJb5H
EIqah6sglOe2QuFO+vq6z1lJkmyfivhxu7oIsELbkU1snHj1qP6cZfsL6aKm4T1Llnw4okgqiXae
vSkSydwCl2myQPBp28af1z8c5WbICxHUFKSWn2z4LN8lBFGxSdnpE2YGDWOa/kERp9rFkyc/myWc
u5okGH78xpDqkpIsQp4AKvd4p9Ibv18Sm9bpPgCaAHVcmgf6yPcCv9ttdpbXo78qSUAL/kvwUEW4
CZUzCV3iQ9qEC5F+Lp9cXeakiRlNParwxKjelcjxItYvYw4gA0Tfcm7HfRsiAZP72g6kSXPH7VqW
8v8ZSJ1CbJ6919ZJI3yz+wVnG8+CIjTcbdmdteuJncyA44qq5lb60Dwyytf+T2LXNh2CeZA532Dk
cc1/2FF/z5lozUp98WazaYyyf6xL6t00GRZm3JTOH4h+vejdI+iDKRAXBQPBn7wvCxXRpxsmL+LB
N0L66Ui//kUGlozQSPJScbPsDuz0hYmBjEuiHrfo5LN83JWQoKOiIsqJQddyeEEVZAsh7mWQv842
1m5K/jeidWrpBexojjd591+I6e+mb3OtxqnlBlBP0eiGVrT/rFJ4/ECm2d8wQMMA0i51Y4NBxmwx
PBdlNLLHz0geHd4MgWTdOw7iES8lzv5g0SalnCaeenUw1KOU/OXgXLOPcvmKZeLvFPwjLYshQOSC
WdvN0K2YBAcSynGmH+rWuWPV24GQsCh4OagiDyyb+c3k+Xk8/6Aqngn65WqA6F075ZPWB+9T081g
/dAIjtQFhrlvxaRZ0IM7GkPZ0Qc//eiLNNvvhF7x0syEevTMtKkBghws8Hi7BhHd51i0H3a/b5vE
qD3wKwsf4JF6Iw1FFzmIXMXBKz55J8gODScNg5UVLbaVoy3S/Q5bdAZQE3jhPCiGQjcVxjvb1svr
DnLFprsFIR7fcJXrGLstqQgncN5emzDObL8A1G6trS/SL49yq8jOlmRz+sJqbLNOwssySdWBWztB
wmUVYfcWqMLSRrpg4kks5vHpCt3weEefNURCFjuQklhlXXRFQFKPH5KVJS/cLi6pGo/fmUHwRtP3
AG4BZ961kgVuh3ai4nkBzDpcx3d3CL4J7wS8S3evmmNHA/MUThkNol2H9Vr5syt61JfpkfuykWwy
8BUApgkWo+EpY8BgLNBqjYCU69D7oyzic9ZiAinMOqDLwuf4YMBLxK+ezETnaQtBJ+CKyyGnYEwP
xL5+2GOYd3eUxiQ6hUZeN01P15j6AU7PNbCCiP214sO95wfEy9SElTErs7ylhbKrVbBS8utIeG5w
23NQU7VBC8lFhDI3WbNTgnskcEMBtpNa3gRsumpnFSRk32HS7RCdz1o31dvpUWgzXzVWqLKIv8MD
6qFVvECetxREzqLxr9nwR7M0cMAvOEzv4CAAhFMn27HZRb4oWSiBt5aBJUFVxYlFQSczN8sshZLw
eBvT1b1ASELeL3w1IOU28/Ctxzp6QaDyq21e9AQty5kSMy4BxWayqwTwWLlxkzfF0noqbXD0AOSQ
FzLKHCd9QkxtU1hFnZDiPrM7Wz9KNZqAkPfGcqsv9BTGasYFLIG2KE+ZnqW6s6/XPz4eEtUFTYgw
NFgwvUld4ujQk1zt0+06Iu8P490vRvOxzya0zDd0oIpVaB8O8ZxRaLz8hUKucWUsp3BnlHnOYtOV
o8KDesAIew25ORviNoesg93/e4GbifxpZzwZL3YdQMy/koxHP1zUoIhCH18jN/xr5CPmniXynGIz
WrC33rrXCJWZMDx9Bl/kqmWmhJltFAnLtCgfXj57klIZY4UtnPsduNUod9PZnSMrZ+u8MYG2RPBN
Q7Dkdg4UDXDvIhN2saqADJbsgrDMWyQ64XjTywYiFFVVMk91kai6mzq/VaYpG3rpoJZ/60HUAtAg
NVCNo56SK+pKufw6bDMA6LnvkyZeeSacjguEHTHMUVsocXsdZq+JHYT/sfYd64xQVaLF0viOUAkd
Ywpwv/TqpsTg7VeXjYsuILWsy9q6QAIwcwRWN/r26Oph4x/AZF/zMXZS8aEKkV6mRPfn7gEOhtkz
TbcMJzf0u7k4sPNB1Pf3xKaKpXAhiCeyYXEclGOv+OpfeiasUeV0h6ANTN4In7aPgcq2godlMM2x
U4V74fZbHcGM1a5EQtdNsl+2wQK1oxDxEScnHLbSDtpmm+h+m3no14uC7QkWoj93ig6B3ECJX4my
nJuMaQob+Op6pg0YMJ6MESKU35IKhFzBfmaR1y/k7k1T4D8ptaF672AicSG4W1wNLwkBLPq+1v0A
kzYG6xlAlFPclhsD1ROm3AZ8vEYg0j2hNu09jmxXxaUD6W10LDMl+XUBjIcfVkP821pnH4KV28JB
N/UL42F9f/sV+W6b4JkPBGeSGB8miT3p70Tc5bl56sy930FROcuEgPa9MkJ3TYYEjnhv408xKnqJ
6r9Fna2I2oNwmqW1ZeMSBEea/ocQjjPAk7rlxU8n3luieFQY1vnVWwCQ3g86jxW1a58xuFv6TiFG
xWAg5ujTAa02i4vkoj8kYSJ8GdWSwH9y5ASl97P7pkzFLz5GKcAkmuPVv3HetgLTnZntueugW51D
nAz9yroYemrXtXjTCfkGKNIIxnlDAoTWlIE80kZ/cpL/bDLCn8fzKHbwXa56zm/VZ5cz3kJFg7Np
aEJlR0vAbfgms1WoWE2w7+QkA/Vizo4egZd9Y7diGq4L1OIXWxuI7ZtkpTXnNT0xKpvGFy/mFGMh
VayvCRDJj6VAk9gHqCHbTU0sjj/NIxl9194HwXr0L6Q5b9L+Ubg/Vxr9MuMo7niaCC7PUUadcLnm
83LyKr3pDCtxJNsczMo0ALkJAvxCO0zfqXNi9hmcx+F2k66aCuSBjpfxSJWASFVDwlYOYoGVaz+U
hovUDqrGn7MJIrt1/6YcYRY8XVdBJsKwvbY2d/zlCNsQCTWTkrRh83IAsa2wKRtJ8UH90vHG5ZRy
Qtju7IR/vNqLi5BEWI49iLPhAFLA83lCukYoQYF7B2onW7vAIZWUHlIMfA2Ia/oR5jaNyaKR4qpa
CZ9IL2KTMQfqosIsR6Hoxd03F9KDsv7xaa1Xbg3JxOl54uYtVMxECRJ8vf8QE9Csmzv304j4KjhS
AbmONuXBpI8hMwHgJbWLD896kpqfKQ1bBsHfYxbC1dphEl2Ium3Hruf5kMgMWnKbShDvkEmZy8yT
5XjP6VMiiKDCsAlmO7YvMY20jF5YDTHocN9E8JsiqGhyvdggMhy7hRVT2GG+q+eGNHWJqgnZmfJR
HWxSTCHEjHxe6JyTUYToDybonQGaNvJeIHqL4t4F86eVi4jdlfe7SHW7+VaGDttqob7B+ceO9McU
6ZALiYWdbMQxXmlaKrC21WGCamj8Yd8cFKmYK5sBxNL72SLJKmW2hvK6SZlL+MhXC4zSzmo6VBXK
57L4seWgub/G9Tmrr4cviNZDpw26iK81QgUi4o+XudppVhYYvBmGYFMUZQFTkMrFAv52oBtlOZy8
jCELYE1HxTBtfMyurttmet/jSx0gFPFgeXtr+PJLBx/uhd0qnk8LJp16Zyt9NzRSRE5LZ9RIGVAO
IUNEYsqRb5fmtgBIfUAQx8UQsfyywKNhGeWOeE9gz2SMDRhobSTFnXGf4QN/dsh3mgz59sUxqLhc
z59GHJWgxrSMNCVBm6qgX9FgWXIfyJ99cUKXDeib6SkeSloIyXZzervWQrAw2ngygnj8Gu5teRmR
sSWZOIQWQyutrdDGgkb80f2OVn7RdgWAx5YL27BlfzGRg9pZaX7tRBuwwkHqCf6XbklaiozmdxJ6
EXsOp1vEYtWcNsbbZApEUUJad1pwk9E42McTEYXQc6eIpiynqgxMuZX4ICH5kWk1UCwX6L311Y7O
QYEFw2r/5dQVZPUl5y0pNTA0ZiNTteZ7IBcG0oT13NOmvQyicE/uKgo9GZX8VCJbOzoEW6p82L/9
XuXhFg9QOOEhtmV+raZWjjmwb2MxiWfg6ZgJDm7JyAmW+EeeoQSNYTTqMrzTOWYT5ijuuW9w3mcc
BhDAPmksIu/zKGQ2A+/I3VKgiADwJEsxZtEbNqcLlKBD8VeZlWltFqY3EcKV+0gSjVfOICXGdu/7
fMfe9gVACSX6UV/IWMUup09EHTtVo/M+D6TyzODhxOynaYAUmTnbkWd9aKXfkYNcAzTMF6Fh0U7t
g/gX5MdMzhyaulDipsQlIXCiKygp9x/B5plarD58IRYHPyREWyIC0WhLeiNnBNnalgKWrx403X0y
wNdWaIz9N2bEsQ10QE2Q78WpT7c6qLWg0Y5n003KqQgZeOXmzQaMJdEiZYnXO1zA62QpaMcIfJTg
32x87u8S5JTlce7RRjslpc+2olvjof2gULd1liQIqcvoLixskAgTwTU56QxwZiMXpyBtikQDtKiL
FauSspaoqs3fu7O3mON3azUxyOHAMz8L5fRfoOTGcsLp4AoSzXK0s54AffrATOkRYJ2Os1o6XaI3
RuU1/hMaf3Il3aUjnxnmvYkRtecmtJ805HOU4bzZ79kgROBJ0BzgDIXnbUscxOY17FjSoUZBFc8z
sbFhIJleJ3QIbalh/f1TNnSzuTSlT3NhZoe1Nfsuicy3ttq+Y8whYdNct2RzpETVtJzJOhtg+smm
hkjuu7DjyfwEguFrekiN6x2VrULRDnSp6lCx/rhyzOnFPL6wqmcvEmXlboVLAFeipUz0XF/wyY6x
5dvwuVayk7OX1yUDIk9RAq7qapR1tRdNZNLKmWyPRHi6l4DrTrephrQJvBalJsBq7qMDTaiYbBL7
D7u9B0G3DLR0aNu4dZ+AFbEUbYUWOZxGuDZGJ/aRO64UMcns9HjmUQ1mnaHgo4cJutgXnoa3EN0n
HZ51dg27wfucdZItZ/wshs1hl9dt96+dgrsT5CTgfZe6A5FHNjADS7H3SA1crKc2HXSiBEMQqVHs
Ay9w2K7X5bxy0/MXfIUduwsoEj2i2LiRYDPdk90HGbiNW/S4E2XgF0gF6PpBMgC4Yiqq9yYbr4Nz
z7FBAED5Q4ZYel5fyaW5zDHvKNovTkZUbNQWLqCEAKerotX6inQ8HpEJjTkygRW7mnJM20vHm/lH
y3eGYfAE17GtVwl4M0JgSBW4c5OMgi0mm9UX7DTJD2hbfnJ1ciaZ94OfpRAwphoyXzjUNDRs9UNW
GLYAR0yNqPH+KlX8BHoSNcvJGynsvyZFLIVpgIg+IaDHtfAfHbPEvxGAN3kQzgIMpTIJZOOn3vm8
it6ROS+w/DCfivQlU/3HFMmKBB1qxmI4Sn+GAQvncWOlsnCBkItyoYm4z0znaz6dgy8+x9UPCAWi
1YlVP+dO7ibrUTiEjAztqIl4hB+emMac9HXUF0oU7WGoVRvfGc+ZkVDaIkA2/otr9Fxri60JGYQO
fPsCxLdm2DpdYv7vdBTlBErnCHHePp/RWIU1npXmkn4AhxWyaB+21hDF43UiWy6ItQ/fH+86YP9d
wbepwuw8S53VgkMgDuSPzfGubDPl+cmxeBvOdKCgN3m/Cg+Dlce8N5a03AA7StR16xIZ0v6vzE+j
q044ejcwijCJcZb6Iwp7Tjzzw5zAEq89ILxNODtKwa5VOOsMDy0ibMibUp303bjdrVYmrW0N3R7a
V5OC5OdVzUyQI0l2tg+GHfGo1bfrXcVT62fsBt4JGAy32OBi7iy4qDmlS+zYfbXEodT39GqPgU+E
KP2rZnp9oqxiDSPBNyLZ+dLKHlmvGj/djdjswFs9HMaOXq2Y/LiIM/S73CKUuHXB1JU4c/C3lG2a
CC+gpswOAuExxUiWCF/zAuQs+g1DvDMi/oUE/od0fixRh3Ku+rsaf5OrFucOInl9S9d1i6Dhc+Zn
dpfgvx/umFexZqC7i6PCC06xt4LkiRsw6GNdcWViur2mRJKDee3k2iC1pwIPZSF2+xx4GR4QO+OK
9jpDKAmityOk+WzsNpzRmAPlc5P2M8GR3kD97Ed0I3klfr/X1Orcx4bzZ4UmmuA+yKzT2DrI+GHz
5umWhpvMxIDti2nEgi4jzxWiZVfZrkPC9jZN6qDFXxkT0bKm+Gc7Dy2s+druVDoVrERdcgcGUoMW
Tf2sVLfdwPq8/fBvFdt4T7/6z1NA1kUqjiVR1WLLBsh+9Zdzgo3ckCYXxZdr7k0ycCSabli3FNeh
D/lrRXZEi+Vs76IBRBIRahSGyqE9RwZdTzFu+JBcl6ZZ0kWwQdrmUovyVV/vQPcwtp5DbOheRFHe
4+tIy8aypZSjRG+AuOoVYnzBoy6LFLVg7Lx38r6Tt864B2k3G+lMU0owjXSAEfrD7L6LuOfFdpXN
GuqJ3t3ApAV6k5yhVXsOe8/xZRIgo81vPfwNeb5pAg+6QWdmETnxc4olr2suBNfLUlWodA/6JilJ
yFE2k83a8LG9RUWT46z0NjNoX6EPyGGAqi/FpYdPdPAK/7S6lXvx2Wp2NUPWzWEAyaV3KMNQX7Ur
epal0SMCMzLfO7dydqwhMxDRx1eoi/6bjpr6CrxjpetPI9N6SPaQA8qg6A+c4ltmpOJ93VGK76zp
aEji0S6ETAH2baXdJeOejGS24JPKX0qHGdqmYk3VKL8u2AqdAaPxNth+IFA8dMXkRbUyMDBNYDx5
mpFpwkJrctwO05w4LaEHF991SGCHu/oFwGFpV/oARA9iu4awRYYPkZkohSA3xycpTOL0ZKGOyfO5
yAMRrwPCC2EtEQDrH8hHVSl3FBWsUHX6WSqMQqVXoq0Mi6yu+bkqCGCAMAmroTQcWbHa9SJ7KoBT
/a0Dv6zKB6woRaruI/VJO4ImBgVb763WYHs9D5JvStbb5OJG/mJUNNCqijrJiWkpjVA+Z1PtiJb+
55whUADxSIwVSQ/Jcv01UVmGdbeXUkQwxrP4RkZ5KWuRcJrDusGswick7HkkkW6ogEaWAsnMdrXV
AKq5kmJDfvtbJZS5NeCE63j7DUu/AruA3d+fYVVCEEmLrtMx0lN4GO+dTn9MyLR2xUlaecAeva+n
v4xUF49hGIX0tGLD4q+E7XyY7SqTrGpHpckR12PVFU7zPhY0Ri+4a35P+lyJXO/8t3C7lkRcRGo0
fTLjzCLLjEK/i0jTJDrsT43yxaKs0eCu9EmfYDOO/IF1702OsYn/yrWA/dTt0WlPsxEzG0H5pIXC
DirM6TOlVFKPAcQfbJW4o3oMF/K4VRoDCk/G8XBpIXc31F4dfDd8IN6MyCpx2jn1/pcRwRs7MMfC
bYHbli72lxSZxcodSbEyv5PKJpDWjU2qa3Zkpmm/CeYHSMa6atzWZO/nLbslb17tzpb6FCncsDOp
oQV98CfkilTDyYPzOAQpPbyUhxCOnZwAVHzhAjCIdBDvSceD8RC1YOq/OwJBs7HeBCz8AsAhX7N+
Gq02D5CFWbWMRPNwJJXwrtyY5ek5Ld+cusB34589w3dq1W3k2Z2QheDb0R7sSDkVJc6YO0qziwwH
epGbPVlelqvx1UobgWsuoTqInf6lvFl4+bYJCmjj3RA5ZMvqFruSixGbEh+pZbeOP0z+TI/Q8s+j
R4pXQS8hcyc9qFR/yUhtSms8QcgRSGST9/BjHEBjXgN/7/9b6qh8hGJvi4UCG3xGwPpQr3nNRPQx
qJZnnb+hpV+YW6hvJ51sMdQJVrTAFv43YNJi8/TxAjTHd7wX1GptWKVXj4oMnYggkh4dDXut3jgp
b5liZuT5l1y/Q4//D4Ohs78+wOJTUWfQFTtdHujs7uoNhZ7Zl28DWHm8Zoab/9n2/Od4nt0AoBMG
PW2YEf1jWG+yoOIHU5zjKvd6rmLswRGegyeGSRd39KyYIo+4zu1iSRO5PEKfEoZLtqimLMHCG+kw
5kOQiNMY52UmoBP6Vp6c+vlshxoufI9w/yGRZ/08CHvUq8Nf+9eQs1JBBcauV46KTM1l/4bNebuC
W08wIPIdIwJ0jcm0WrbJ0wGiyjsTS/uYX+x1rlk8RzfSgdC/1/AuWqEYZWeGdct/Q6DJr/LJCbgc
hA/Yz2yxsLSK8+gbs9tn79NTwk8s+ylBiMk6nqwP9YBqNT3m25nGRIpl5+lkAi/UDBOB321K6vxY
kHzcoiX/l7vzmqhJ2hgztDF9QIwB/xSz0XDLcdRqO54OjEpi7V1hSos4yXNLwt7pNwvSViSOA0GX
lwIv+xuKNB1H273/d3JekrOEv+bF09K8CFEhBFhbQ+QRpWFkxVsTE2uLY+dtVORBRBsbuBcF1U3/
bRnsrBPwOtCO1I3pE+XNur/Brnabzf72HTWquUv996KuOmvtnxlfRjqsFZcNLb+FoomW8hHF1UNU
HIigZjp/Y6BKefGBQIk5GkurCyU9doYByr0t1tpaoM/twjPpSvtrqi1MZGgQEyfg+nT0aCFyCdhU
Biu01ojx+eo8S6p9OEj2pBzGogseL6qNogPaOLBC+rUU6yWucY5BxOr7Vs4VTh/qd3T+wecHV/uE
yex1IlVOeh2mSHm/pQKotFldjyo+A2v0xqXsE/pf2faamkKwVpJhfm7e+cHWOWC1Mxpq8qiknCOz
/1TMNvHwmmd9PhvukxX0F61krQdSiJEilqZa87Qeb4bwQbkvzVh3PlE4CsfUI7piaDHvNz9tdQmn
4tqR4Z7xtnTdZB7LZI7MV0oVDcebYTg/0buYaXBqTC8+U/Ib90nU16/B6YwreytRtbCXw1okBMGi
DRwEzjKKPQ26l2dtcS1gMKEc3kIgh5SpjTWLuabhQ2ZmHGc1QdXYTgcUzyCj5KQ6xQHCp6MiMULq
0u9FmHMGckuYhhJayKAMtCp5Lcbz41yOaKQk1YbzFjYiM3nj0Qc99jB4gZWINd7LWbj6Bk0q4c60
zrNcnnoRTHwkQr5fTA5F80MS0PRpP7ZREiXnroRgcnboS5dyhTQQGGN/+zy5Vd8m4HDE4wLgkCGx
L+2y2PVB5rdcjh/NrF2niNkQmuZlXgcXOHmjekR5zXFrpT8oXGkeUWxfZIa5GKqmBV5kPnjmvrrx
B72i4a7Ccy+EqT5UVI00N8mvLo+88sgIYLfTT8rGgqoqratQneoQIkcQl0z+Iq/eP8HpzH7IT6G4
Xej6r3OQvduWcxBx6GZRFjc/QlTIBz74gAp89Gs/QfRbCW6mhgNtZHDXSAw1TMT7NztFk6o9wtfb
p9iFWWWOCthqchkIwHIo6ngTTCHZgLF5X/74W+dkE0RsKIpAG+aa/2yyp24LrPAoAqBlhxHiWnFF
nXR3mGJGO82IWm1NNxYSwSTVlc+eT+0UZBGodMrLP72cOXRn4jJUCqqyiVYQHf2EoOTME7vKPNZP
TyXzVnVUzZTyRFaKQIQbSkrH6XLC+BP+wUfGtZO5Z46QlLPWaCwph8h2jjk5eT91bC6X4kSlMatF
fZRqodiuiyvELdNp/tuh6ESFoi0cEyriDuTzFOVT75R08y4tDiBe0n6SHdYI4fYX+rB47vuVPjKx
HtdKHmHVW0p6zGbtcKEdbz6jLhYKYzQgv9DP4J0ONayyOJExZwFOtN0uRzh82Ofps5CoLHmzO1DY
cXFJnBO/4Rhc0SBWMZ8uNaSId2lXhhRNLlyAe4OrZWeVWbXe14vDMUgtyBUcvVRnhPsPv1i0JVRs
OMro0Rr/CJvUPnuqlkizLp1+xMKpbxZSi8V7n99xTGxpZHiyv8uLswAFwgsVPcSY+/xQtsLv+kDz
A0Rfz6tfL/yAQpPhEsq69NH1orS37uKWgq7ff7i8vvPz/svm9j/H89NGp02uu8DD1iasWGG1rcN4
3yuLyc6emR0Oz+yMExu1O//ProkfGMpqlB5Nt09an0vrtsKfT5r7ybt2LzIlStslNUWvwlRAtFvU
zDE55+g3+jctyH2G63aK1M1lODDwBY211eNuV5bDejHlWg+KteqYUMh2H2YLL4PhruLXoc+FLjMV
Bmk8hq0BRPtLMC2cwsgOqrwUG10zD9aB+Mzz0iI6lKGnp8xxkPnuCpueOpD+sHnve2aIwg2bwmOZ
bv5GxIZMsFYJBEm5v32PLjMtE0tLFIFzr9avbcmDP5WUG8oSDfaNGp9a7cOTNP948dIckAhf64pB
mBU/mBaNeHv9gdq5QS7YZ+Q8Zlg+AXFKCXcbro+COL9ryV2eEPmxrSAg0VzVZPpT8Nyhs9ykjWqA
YLK9ecJdr7S8Xk9s398r8fUxGPcZWV6/vSegwlaSY4trfWW1U1NGcHRLPnEvPMN5pDMb9keeApP1
/2C0OdpXbQuY+ozv7oHLAlv2v7Zx4HUPiDNYbLKuszliQkiiLC3lTbQnZfLgOtNwaHee3P+b/IK1
5lIi1TYWSThwB9Rz4u3HR53/BU/y/VgBQTp1jNQxoz3ME+D7jQ/7dwWOqDP1aRHrOZdWbnpkGAsB
3v/jvHyc1/qrWP35z+QZ7Ek31dxxISBB3QBE7L8eEinIdl4aFI/fHW74cRSInDlPh2YBgmJrtQR7
53bvn7lOwffXrAuOH2ykqWrBTGBLnkqQBNP5Y4IM1CAM1guhRLYGl6IzWuph5zJyTSMT915Wa6P9
fDReSan+gAvo4cjtq6NvVeC5B0O5R5YY/jEmedRkPA2S/akaV7Ts/UyA956lvwzUDWyTT9fekE37
CIBQFkSoc4g8cdGp3c0J5XFRIctXqNAgGOKllFajEgL3zSZ471qFuOrnk1EWn36RPrrwenqURma0
VvRpsqr3eTCnI47R97Jl/QpCxb7px4FWAhNmu3PweeZyiNbAQL580s9KYTZFX+Y1EGqJ4wbWMPM+
7yTpzJwCPec+h3vboz9l+kifULTtQuoTWgF8yKWRwwbpLxUgo3MncJLx4rWdvwMREbCj1LDh+LbY
dK1oEc8KmQl6dvpeO8k0JaPWaUmpdBY7/VDr7A7KUfc88zEVV5UVgvQ/nk+N9Skc/KLi9PI/6num
gvy1Yalts2W3BY6b+hjFLGsrurzp9+9LxBaavq6YafffiycxyNKvTinj+P/t9sZaCUcI4G7RDIF1
yGf4XBp/kHq/dio8dFoPYnTuHV8R6KANOX6Jwc+u/wmsRhCyuCeBKiEs5Ey7UTOZDgJIEcq7tIgO
c7VljNctlENnZ9ucCyJFsQHgqV8NLlOiDxgEjpG0b6gNgWLWGZ7b+XKYUctpB1bxm2+YxK1i6vGH
AQoZaDaE6jviVAum0HpGP02vNpDmdo/PgTm4tJlBzoDYODHp9LXmQTy33S/HFq8x7YjDMWXs3xox
Jz47MqCfKzBvAYKUCSIr/0qwP4W9MMwodUk56YXQE4R7zkyPqonOSyeaw6ERvvFGJjAG0Kbyb65o
yH3JAozYb6n92RNKWdkNS+RAPYsL90RKPmPwZxEosr7uJT/ZwRL/ZGZUiVJtt7BSzW1NdAxAcWjM
icsHLIaDIYKkl6boJV4GLaUDF2ykvudcyznWVH3IBmA0LeoQit8zsMzTzN32chnJ7aOqAfyRMQak
FmbJUBMmg3abcbCBVpI08sXd0eVX3qhncG/TAkOhMt2j6jxLRfOeyoMLDARcATgCtfEFrNT1R+p7
whgeIEimMjDtlW/XpsE456MMijxIBm6jviyiKFgqCfY8D5DC16SpXOS63+oY66kEcQq/RXJhyXQp
Ksm5YXYZuj9NMUPHKphGjwQ/uGG4ep1DWYCtim9vmfrEWRB7tOpPxtCCxGP1Ma5Pue2xNJnA+p+3
1FyZAOSgmHppPVH6fqb8VrewiCvdcMvlR28D9qeyoin9jsSXILXSjr/WC6UP3tr48wJQF8ee1jKh
/G9b/CZUKZwyOQx/GDsVtOzqNKwPjlo9YsBgxhtcmvSNaCN5WvhZeN3zEdTrtfJwY4z1ExnUB0ui
PYO9KBhPnUK64lkyeQg3rquiaD9U5DOTstYfkmdD5sX2pKkaB4hp2SLwQIwVFMy/PlJeMNTRzfJN
SUGmrfVUPPiflJ5U8J1/IcgiZ6lK25LmzTOkhiW+JOF0CboCVMrF2KjcUQQVNbCpVBypJA5PUi6Y
a5Lk+DPvWVJcXlHJ/CbJ9b28Aba77wYx+/Uyzs8InqQD6VWY1QLzcArqo8b50D7yOC7ubWshp958
Llif93/IL02E3QjA2H9b3sYRsA8bt+0KUB0lwcvNb8hE1INnF4EhnMxmZMy3upxNivVYrSVqSu70
ZYMYhC/46OINF/ByRA3PRd/edOdK6LGjDZQumYDMPnt/boVDmJ+PUL57eDo/SoWJ3IjUADR6fHb1
/mWMNf02H5gCRcytzdHlX1ExJvwB+UJe87HVMgJ0j1EML8WewRutSaCF0aMZN9YO1dgp2emM+eEF
ZIgYbclmEy7GdT9xTPmhDi0vUzpng8x4LZCDbNUNQWroEJ1uRM8OalbI773ReIi9kcVNLZ0m6f8F
fh+SKJVJLL5kRNfppHmPi8+UlVoH4n0XXE7NW/92/dY6Yv8yhCr5/YkjxF3u5zBDuXKVGcazTdpT
Dcu8iZsQY2bfX1ZimIqrAWGR4Y6SPlJojNAOFhVCD6Jv6SDRda75fE6Xfabr9ZhA7DzE4UxfInfH
kUkJwk+GiggAZp3G7slCXet51kLrp5Bb0Zfu7RD5WFpzbU4Nwxg9CwK13Zh6Dx/Y7LnBw3pRv/Uu
caq2XLsneFwjot/niiOOwSJHmRyy6frov+rbJzZLe63xV+40CQkP+Dx+8jQAd/grFKRvuD6jrZTw
v1MaJpLFi0dU3evRflNzyBMb/ZljcyykSJT6l9TbUSfmRyh/omC4peXRJtTQZ0w+bnhj+aRY/pO5
zzmPv3VM+whUEsP0Vzq735upLu1B+kchfIgRuOY6nb8B4PVy0W9GfiNjaL9pgXSLF3x9gKeiA4kd
4I1/FQmuUkx/FIyfh7oJbN0eAXm6vytouxNCqCUyr3k75snlAbTzLh5JkIK6RQHJOOCji1jNmdF3
FfHrMh6LrFU4Kz96lgx4P33oMerdd4/jCyH9nQg9vb+NyzuQ8ByRMBcMXVye3zUNCjf7z6NHwoTC
WChK5wv1UWFlXUBEuxTcmlo1q/ZPYRD21l1RnrI01LTLwsfFSUUCUc7YQtAw+t8XdPMLR+5sQcdP
TXKjOSx0qrya+0oxHFQ1cV6Yx2FIWXlRes35in/DI+1nyhnnwlkBYgYjDizi8pF0Ztmo9km4AgUq
VPqJG0dPVwLPmqRmS5gbsh83oKYODr+coZwG+1JWoWUP3JcgxiP0poacnmRo/+BDkqYmtGjRZGu3
Adih4DXCi59rjqkLAMYRh4aMFD0WJXfEqlJiq+w0+7aHfX0/3KFqfq5AvmvktYQhAyo9j4SDluqx
VP8AN5p8h54POxBQPxjGi1B5DfW4PyMCevW+qhwSvRnbndyvjTSFA11DtzRl24spGIV//eibtc+1
ynv3mW9nlWONVTxTocYzdgwLsbDCvY3iuto9hKG2exSpga49Jn7JlDL6cIOnpmwyQb25DSoo/M4u
v7oD90jVrsxinNjF5yRB7lfS3TwmrZouf5okQlX7IXLBu1MoAcFAMtIAYQeN67eBx5s+Wdyq46k+
Noex2LrsyzsM6Hpx4YqF/zfStl95nQT8ORyOJl4qccsV5qBshvIBK0vW/XHjU75kmqP5nzj6vKc6
f/WJSCtkIMwG3mlIYQBRiu+8eb22EQCNLiHQpR3bxED+FdAl3XVpsiPII1zV2lcYLfg15dJrXTqm
1LkyE+j8RZCznn+JCEIyod1QX+ytL7Q89ZC3rFpMD01kxQmu5Cjs4veczZM6ij/kmNMf/LdW7v6c
/MeAVmf/CykVVKwLTdBWT0DkgHC7vW+qVQnevA7sKGi6PnApXPakukfiDDXFNKpRiy7Kh90W6c50
0J+2bpEHbGGAyo7jTuId68RpvLE9N6dGy2q0qCMEI5z4kCYHJ6YLYNuiQmrVMsd1w87JROobTGr3
jrnOEwiB/R5wEGBSq2y9SVBHDDYvcAoYIx9mFAL23rx5K1xqK7qCmysUbsyCUSEwdYs09b7JjDuc
ZUPy2Ic8ri+VXiPuxEMzIpPtHkbRTvXJVrYKF5vIUzF2afq44Hazim6+hQQFfF8Vh7aQF/kc2IVV
fv3xNgMVb5pdb9uWr2hTiHM8ZmKipXNpgt/taunnMOggR3sitJK0P5QNcbSicJM1nXnwH4RKh17k
NW4zaCpieP6SvyRS4OfGy0TGWn/RDR9LOyZAX1ROGS+6Kuq/JCBQLFAHDbs7gntPjYu5K7ptoM+k
qHHBR3r6UXaf2CzHqgAsMgnxYmdHHwl3YcP2JwLr1DdVwdt1vA07IJQSEo8hHi5xZwYLX1l6zl1E
Wc/eR/NjElfVT4+DfKEBP3Sfewgb5I7xgHvcDMuTGuYZcv7LitNAXh36F/phine5ym70w7cRz9Lz
zg/JUDd2OwJYpJPnJkH8MIjFsF0ZeKuQqcDjGKHjqvIkhFCyW1Fz598PjT9Uf0P2B15J1OpRzAvf
/TCwyISaQR/U+boXGPXPiUaQU4E3fKbc3vqplJuiT2p6Gl2WcvOFzDjkOKYQy5VJ9bLes/XX6Z7P
1aWahSkRkvGxn+FdIp2UPmf3SZwkVQmSwIa+uVx6u8tqjgHTvGXTS0s66EMSxVYuauMAfvj3OIla
REn/kp9Jaoqlhxk3XB3JDjjAAahYmzT/LruoK+eM9fQap7BMSuNqFxsruA8FBOC45kQrcnk78HU/
F0Y3uW4W3I/L7ocXejJthyoKsuUbZgxgbBWZ7YYiEgUVUoKlhWNY1EyMUKx4H3IFYKqW5rAsoiKx
9TUhpTqrqfhGxsWgVENio8DXvvKwtskJw0uhRMdr/POk820FKGEzVd1mgvrsdsiN4JQNZWzFCFLM
esvQ/fp8oKnTeV/jQ1MJbfiRZTaPhbuyoM75Kv41V7oTSpkXtNQFHKWoA1lMAWW5RfDj1MkHrMjB
7Q/9sd0ib40pLJg/WMPrxbRgL5uGszbPqmDamu1dpjDXARxth0G2VyXGzw619XgirNlva80ZbGq/
24EdVYZTtv3ra7vjMovkywHU4nDGCNiMXFCzdYCB6egmyYs4BdsHBHigb+C3KnbQasPW+XgxzCNk
hksjddOiXpliMKehO4qZNbdXN6C8508GsUtNEE5zInfw6zeywJ/ix9yPmG2ZnRaCUQbGDqYnZ6fg
RB2EdNAhSNyLRNpsvhwyBu01Ad16itlycMaG9gvRZjbR8M7WYaAcjIP+fX43qZFgH8dojEEwYk8V
OJP0nOcBmtnp9pWBqmD/O5MYi44liuPeXH7Z46/5Kvg5GgxAsftY+KCKZ9c1mzRJAxWEnLWLDmxo
bBQIo2CkGH2Y0LH5sqFjwgAPRkAzW7vSobxkPES40WTItgQKMlu2n5n2cvuYxD8Bi8g/Z5hTFsBb
jao13vS9VEOEktjGUjXSFAefHYFB1weASFWQ4aSvodlmd3n5bMZOe/CHHu9+ixR5pNaq8ymwR+Bm
Y//QtxkO09+WRoBpBLDSggZTOYYBeta98vCMJ4KrjtpSDO881TM+zCeCZS5C9B18LNW25ZREF3+2
d8sNZb7Xvu7aMSsqH4go0o4kRtoqKzhlhT7YLoOoj7qId/Qk+yGxnn40aH0d8dXd+k6KaacZlRpK
IRcwS2NMdxcgGb4tTvk5V5jBUcDkVTPT7niBKnQCUktmyYYAyjWhdx9oxWiJ7LbLYUvQ9j++R+rp
WseQXFGCr9awSK1frmfA8iazfwyQ4WhL3Y5ENATwBV7abW6IknWep/50rsOsQW7aMtfqdhuSM1Kw
/fTCW5H4fJbcEiGQRuXDOXWWXKizdoKX6LEhagn6ap9k1MNvaOcjkH6TOxGaL264GNkfe+Z8q4Um
iKZRHfMufSLIx63isRoHLpemFCK4WpuPPH85S1krEF9o9+lM2BQDpCw6t71Row+JxUes5i86O4fv
Ko1h5asRPfnEVvLnfJW4fFNtXBK/Fa0eZSO6Mz0NetEJ72zBop005sDsHy/zBTW7a7HNisezrh7D
ITdbefM5MWf8Xbv8ewrfL9WKCt0CNEtM0Ah/gdqOgCBW6Im1qPUqjbQmP/YDaIe0PutEIZvvQyUi
AlObbBJn94nVBLW+0vN9PPAOIEnX9qT09fkYzfz4uj0HxD9O+Ct+dFc3ZiKbFLeEmpgkND0uitFM
KQ2Xyo8RAHPTpKQ+Z/5MudgdANLW+IQC1XIFpA8n7J0YTQwwBmmmWxVp4k/PYKpnPA55JLlvhM82
hTphIkEipnaK7w4a22H1/4z6ptIapYxne6RurfP6+wJ7GQBY5ecJ8qeB3U9IoMHmMTLTPPY6YFE9
+OZ9Z+u4yy9sgHnGK6fE5TjkG6WQ8+m+IUQL4/VoX8prwGaiPhAw0R53HdCp0fr6qYeOPse7bhRE
soKYoQOt3Qr5hsrjEVlys1Qc4uV5ECk5KpWMAIuzGoOiFGbUyavsLC0N6MhyP7lwBad7TFucnD2K
vQmI2Ca8i7zg6HEx9lEC3okoLvTU9hOreXVN/01B5sFg0oj6bZSUJ9cgEuL5vvF/GO/uomsVye2E
UQsbq2AYvau80UmsurEwQaXG0tJE8UCixBDmIYXlb5i/KwvJMpo6evENHCPYJiOIkitVjyyqsOK0
5jDk3Bw0uJunVB+eespjonMLobxUMhbp5Eo/yl/hsoWfZD+Lu6Ij/bp3V93VQwncjcMpJVk+hOY2
yMeJ/eh7OsZ5ebx9vylJ95/adQtDQ01t9Ms+vbLO7EjTOKa1DSd4LQuljH66L/wjb6raYGeNWKbf
2zCxyUhZfFqFRXp0V++Hsa8sFF/n9gKFgsSisT20MkH1Z5tnhjgeU8uRPz5n205K8C8s5hruMfBm
acGUWF+R0qnoxcIQUjy3koGA5kvrAr2AfwmXqTDtj2ZaHngim+WXZxQTycXFmWNiV67b2rY8OGj+
XwNJwa5eb/zahEJ0pD1/Xv5uNmm18OJgdkeEU6qCkcrX7wvwt+SlZbkzaMFHYRVLPAZUkg2yJhJp
3KrKN2yMhUL3gmM2cGIJXmx84c9hFJ25dnlNY+YkktZexKqPrc05O+crWTj2CHGDRdPyg/PdDawH
AEpeVxDoKb4vld/wm8S6s9Zo8EbcvkBG6layQFMzpFBtirm6kCADASxg/CKjg/y52idSXx/8q+IG
03LbQtmSCb/C9Og9wlreh7jhN0R0i1hRtJVw0V4PW9pDiQfY9XP1i7dPdn4J7gS1S9+xs7bIQJLA
VcJn57F1d4NISqfH3yvuXIpXmMGx/eZA0WXHo4xVI8y1HqiXVY5VQRCt+9LJCr69Hc35E143Mjdj
vSQWplsjoONwiApK8efdA7nDTLrDTLReUhptuH0608tI97vNalm+fJdM0thU3LE7fn+vjzLuBcDF
yR5L4MgY3U8RJUgMlfJ1YIaZwSP0dwFxuLOV3Xg9SMxnu0/fNoDS/7WGNl86D1FeplX+8dJ7VkSQ
uMRzNhZwFvD964skWyiEUPdQZpN4W+ZeKjRQQTYrWLxFwL16m5F2qcIDXnocr/QreFq9xw8XXdlA
UdOSUIVpZfpIFTinR04t1PkI6fkypmcUF3jJEKyYAiFNsUz1SWFQM/6XGsBkr1MZjtTjffCgmQTs
WYXhAra4aIrSEIa16+SpO9oSI7EjotRYohzKisg3N3FzZJDGloLpOBz/+pkgmnN6DiTxoIwsv2OG
PUQe+Ki6rGTLRMsDwB0kaHGp7+y1TYHOMkAS9coZ2gfeDazO7k0g16wOylcr+NjB5idt4XH0Wr3Z
urMAD47oL3vtWO0n8ooWS0pdU//02VaRp9D7fI1H1d1Ga3ixuG4Zd7hKaSCZqSMlh55kofbtVsZM
tsXRTSR3x0O1xPXjIQBSWmJZ6J3zHJ8XU5Jz53fAs2KFbQ8fuDbBhtIwxICx916zkjArXmVbSH15
taa+jxF/Vq/+dbwAf+hDHEiNSlOBYN0Cf4BbDkkz9PGXtiUS5ybncPrvGn8/O6mIJuzpXAqtBiKs
CCv/4bzDIphQnsdfNAZ3M7yMmqlJOwgfWOmZfHjg4jKJG8iLptu+UA+K+5p7Fveco0tVa+7iMaZl
MLrjhy4EZcT94czvwVVCtlomv4Ph6d0SkFxnK3JL/MpwtDcpVWMOCWI0yq78zBxbs+aKqosUMVc/
OEyy/g4cwsiMlk3EVwMq8+lpC63UHfYJEgqsxoMU57q1jFQIpFXZLh3zfbUP1fc4QuZi7qt6uw3Y
KYU1yvl0+jCRoJhuAbZhQTpE2CwQ+jKNOVFr6B2UELBcvwC/1Mj7GNE0FjCKO6+3fXYjf3/ZlAFi
kheXKrJpukeqOxxKrLrYYnPtbZ5LQsrJgUFNzcCOax9CIfPqHq6BIZCaBST+I31Yz1kWU+XT4Llt
QmXGGXP83kqK7OeQN3OMJfQsWEA8wVt6fkoU2rQnMDU3gt5CK+m0bwwQrNZUf8G5+5iN3LYlYKKz
ClrS18JgWX9w0Pua38JaP5vpN9kMtL2RIh1alCuYQ3gl24Kp/RL3tfadXUyJ2BoNnxVgOQHf4wSQ
JAjVaoBjehQZEab9Cu8fkjLhDFlxOv6jmU7EShKab4XRDWAkTPmK2xG6u16N6ql+E9+pi5GwLwCS
FSH0piQr3qda72bkzeY9WQwFSfzriWXmkx1GSQ/MB2CvUBpSATxzsjIIB8WK7UOikQrBXznihonv
wXDtCfMGmevhcTvwcyQ6mIoUKc1ijgBv+r+YS0Hef3tM+XhDXZTk35jFMbeso5JhnS9cXQTmhk5P
e91cLv08bAu571GlNinSDhKRvPuA+zATwFWoignPl4gPXeUFP2iH5uuzQuMT3UjplRj+mdueo0jn
SI3DzFqvrj3ojPtdYZkji8egx2k3npC4qdNcQv6BXAYAQtE1BKolqRSbTYLRxpSUgR+tgnLdhhsY
mhbOkQ0/HoT6A6MJkKQvsrdvE0w/X0yflvooF/QPdjfU8+Et+Mf698hBa27Yud+HpJunKCSpVFAB
pB+soo/EvJ32TLWqTzNkTOQrD6LyAZ3R07R5hXjnA39YLL6DXrptIWowQJCwyZbMDvvfxj36FFWS
GrFCllLwGktjzLxdQl0Als/+I+zyHPxXtfi4JFV65HIaps3vqvPLOIWKLoo36AoZ93qKE/CccgaT
lK4Kt/LvjT6C7BIdNK1oiU71BX+hoq71DdaNefxiPVLj8w8iblqAr4+qxzFlXA8y0xxFxYRdHSSd
+2QR5V0ma+E95Z9qifq+Ec46eTOhYjEFCvAmS1Zbo8Li1Kx+TUkibCNX5cHomxR67TaDOLHSbcZD
dwmpbuqumMpVU3BBO3dhMhV4cN/1boaoTB6K4CZnzCaX/pDmG60IUg8OnrW8m4uAq5T5t56ENJoF
GfK7gPYW0lZVb0IH0SlWnmOt3LxWhXLfuBis2OxrpKXTTs4HZ2X2KIG4XhzhkzRbrtfh9tMRX/ch
NjCz+ZIQ4u3bpreUoEeU1jDU3z/rj2VMf5w1y0YxtcmTjxFn/J4QA8UXxeZo98e7/LsRgLtKUmpr
zYFf9tHqq0RjhmyyXL0c3Y9u/Hcu93kinJNc2vyv61bXRX+aU4GVkxl1aZptrTHxe50f4CBDfZow
R0Iyb2vh7mP31N7EJbNw9JMbaKeXyjPbNszQxVMQChWMPWdDshc0EsNy9+7GTCt8+rrevOsMXJB0
k4SbNtMGkDEe+AwTuwYF3Hc0SgEfIrBm7f5Ecvgz6LZuaZY0heSnfr8qUb4oGN+xSd9WKu0BgtQt
KtshJlaJMu9z6Y1kx8JMvypGWBusjoIdYCUZvaooOG/ZnOMALpaimPwuIMQhEioal/F5aTwo7TrR
95agHA5ffEsbBhsMs/ooRUDuCJIgKWU0ygIqDqbucr+7DVIJ1wX/c0nR3pMkbwt8jJTKH9CvpTcG
WHSMHnnLJB2J5lul0aoE3MxOKgfNDh2ivUo/jiScD44lcmhI/kUOrGfQN+ih/uS6woE5cmWcOp5p
rpKQkN7O6wWV3zovG2zvCL3Gh5iiBirCcIurdNoU1U9BUjRG2pfgNLNQ6M2zVHty4Sc/hq9bq0Kg
3ve8Bsgp0T+ZBXm4sDLlVpH4OQi3MczCbR4y8PaqNiDs7tRuxNU187gpCbaIaD1NaI/97EUDxu5w
u9jBjM/bSO5PooQ5bNmqxM0g3/mjxidjQS5zQyKKaCXmJLo7VVVlZYuM/Xcwr4vxUPqxAMIy2o4D
IXuZR0grDRJ3Ux58a08SSlbKe0DK184LCWRHQtSsS385+Fqn2f+8dRf/6p6csW4N/vMmoAT0jYeC
dK/L85OMHsG4D996W0r3nuWICSzsr6Ww8vyLc85ueW71/SlFqje2Htp/O67fWlL+91puxJkO7TfS
JAwmjZlqG3EyuBbel2X68qxULGB7+Uaw7gx2K/1ox0NcqFyv5O+ZfV3zcvnWyTp1Sa+oy5IJX5en
fhec97O/1kK3pwAVmI2NIOEZ4Oz/3ES6sQ4A6DUkZ1ZXnUTpVeuuXhNH9PY8IMQrLSnW+nK8gYS9
3JfiwvEryWBlmt3MBjpBpSBoB8xErdo/G07XUgMFZ+Nl/qG7BKvM8J3cltbLZd0pGHnt0skUq8Q1
Phn9NaY7ruHsg+wHCpCIHWDh9EtquWLrYi5vBHvGUkv3uLoIYar8gewQihUSkRHy6iH+dGmZkcL5
Ggwh9zEOixLXcrJXnrtpjxE2Usc4Rz5RB27SGlQjc9sTKQI1ILkT9m1unO/VLFZHUO4TKVAARu9m
/Yl4PPHALzB+9DUhAzvLLB0k7qwAJEliz36vVtlxVP6+E3cWw+ew7g1oJ7JXt2fpih8IKldUODjU
vqQcb6pQNl08vakBgogZYcg/u8G9H8Lod+n2gaeFmUchrAX2oHBYsSjwsbdDOKy/+d912z+WKHy4
2QKGsQgHzITq5BSKNcw1apOohkCWeyNfA46hIQTk8sQNk0doWY89u/WFmb7fAOK7z2O3fEXUkGLz
sYQr3J9OlPxOm27fR8aEZmC4sNfT9KnuPjCeutretCrGvSa3RSCF95/H1E5VTZJFWjcGOqGDZp3d
53IpYmAMb8J/EZ9auVyhheuD4E1Cc1pfqKtwa210GsO0IwABb/+iOMZDkt0cDWWc9Fe4EvNKHUmu
wH8XCFxv6DK7Ku/DHjHm0HW8pYyITyCB4fRoN0PWHVbiEyOuGLF0b5OXqwCIwBF5tUmny/p9/ITR
HuSEFsanBcGC7SOwxt/E+msZow5oNCt1uOmqGATZBFasjb7OOLzugEOvkb9c8AwXvnl6AH6GJW28
DaG+AnsMIAj9CFb27s4JDy0quSXLbNYOKj1anXrDq8YI8YOk8nq9K48YNLhAzM6mawRtUueUUUai
FpyR/dRV3EY+oZhb1v8H1CarJW+OZMTL9tzoYod4kHL0vhITNaYvHlVqWC7AZ9ZgmzRJGArb9gp8
flwkWNxnSSiyix9aZ4iRuvgQfgNzkAwooQaQIlXFk6pKRMwk2TtJcIW9vq6YLQim+f4Rh0Pdv5LY
5hPg8ZXAddifmM/EPyBS9eyjNzHxMs3vRItiD9s+oeOD41QAtrVRea06sUA5Q0Y9Mh7g8vldlJdm
PGsWLH/Fba6bsAWlNT+HCFKyHEBVkx0u888tLlSY6T7aPoMnx2AGC+xwmVcUs1UOr0/AnryXnZ6L
RjxdksyzFR/pydkwo+5nKvn5xvWy2AjAZgqXE06x4GNFl/CmycRQ6RW7kEFDT4x+/ngMflq7zKWy
D6+FwXbga2ilszfd3ywd0wh4tQ0cPTwL17ukY4fla1cjneXEpgM+TAIBfwLsZg1+DaNkcjlqZOlD
xBhpcFdC8z5o0mNDxy2+pKq11FhdLM2x+nBtUs/ZbVQ9sszEeBTX8m48OqRFwAlBX9BnvSF/bsHh
M7JGK9M7k/CqPmbsMgubdiKhkbwBLsE1eOShOVr2LZ00uQ1bor8Sy+Kk7udIUG3+rWrlUxwApLPS
agOQgf6wEvFyihqwDt48MNMhZEV1r71xQeup6UZFLlRymLybpJNaytpmVE9y7JGYWkw0hvoewtS6
rLk1aI/CeTAoEsuV/vo7L2dwoOY5/WGWb701/u2jlypdFTnVZ8cNqU9srC9DJEaVgT7ldUeEPjWk
fT5ZGI1hAGZrVpESU9Ju2Iiwqjepcb2BvJBX2LZjy5Q49fu0by64zhcRr9D9ilFvZ3YLCvgsFaij
24Gk1fNCJn0BLdBkl5ISc1VzJZQ7Ywg9IjLGPQnwISA++LUzS+j/g9rzLBIN6F7ltHn7gvIPw43q
DZveEGC3yLvvkkPBFaIpfe2omYGX9P3wmLiQulhF1HB0vnL6bllQdw6MxxPfFyQ8dxMo5KHgFcvI
zP29bcAUif69aLuoWS7/c8YPT1JvgGspQjSJ+xdoapxCj8vailEun9juJUg+cgoaNlTTJwNj9YWR
94MXu5s+wl6c5ghlMl41i9+Du//q1OcH5a0KK/IkKXebTpzz3HxYCsaWy5+Hfr2mpzJGzsu5yKwn
3HNwiGF73/xCzXooWoJwyAm0H54AuCG/u7NqjKiCUV9P8hotH2wmeR8xQ5Ky3H6s3Ka8Y9+xK67u
jmM4NAGgUY5OD5Dh1gYsS4iFZLwlOzw7+c0NTQG8QrlttBbOuRQg/RLnAqmMmrd3LVzIaJqz8oMr
WfoA8uYE3DQqOsfGWx9N+wz94hycW0Xb/2h23gkGVWGmwsQY9XZzwi3Ukp4oC/QqyZuGbXoAr4Zx
s15CX44llmtkzJA/0H7J2WD+NaI2NUuTwWN5brzG/2ZuqPB5hPpxB+ph0atH3w/PfYowMdC6oH5r
i+YBG5UNupiHBeXDttjj/TSc2AWy+dl5Hnfw2gz5GR3/jq0nJxLcI9NTQ6bLKbE2YV9fgntq45vv
KgVCWKr/6Hgx2jwlCaMK9j0VhG0vKT+irnVVBGKbQ9w8kGc57royIxrzfIOMOiosKo3cABKk1FhC
wFe6pqhS3WchgciP1wG5aruw8neEMnkVViqOd3D45PiKlzKvEKgBxmsAt65i+OGyr04uD2mEmNkv
mqYluCCNc+fxn+V0uwvoJ3bOZy2nC9nQJIvnPXb8MLIbbo+XyN9ltZe0tw1KpWgtKY/B0e4ZTw4/
pNn5r7ZJooh2otXVPjU1wxwvnMagYQjky4jP0Ifd+M85pzdWS36jLzX2xbx66XA/CJR7RI74ukSI
+blVXAhMGIC4AWfzrEkx/7Sc+gwsBHxKLgEYJ2MpTuwnPX92w9gEqMH2xaeqgd05Pwoo4tm4or3u
5OIHvcxGW7OiB9PHLqbRrTPeZ/1W7fl+aI7BFte4KcBTQ8y27KEMvoinUJmaOLCv6fv/IqqjEBoR
mp4V1wk2/zFu3pwpzwamrIo2/ilgiRXBQbg5Uf1JpAP1i9LRsfBHkJij7WcrvU8OdOk8XImT+scf
CDl5m8ZrBSR1QWJCZ6q4rVckYaDNT5NNx5tZAN86UgyQQKaql8FEjBuTMWynSTzyIvYbmNRI9LNd
ePDODb/pBu7aiadbcMJPXy8jONYRWtN0IJC1ngeuBJGLSCwIqFl53PzhTFt6R7a4E/BSWYn2pPML
WfQwMCetOpk3cSIcrjpZjAUOWXGad92YymN7h8CtrrlM+lC3zaktxHlr3BeIJ4++oJxU8x+Hxfuc
iOVTbwPhRjkZw/qXBRY//EXOMMIDKj2MDH05rDHjU8EzfGErbRjJyNrKSeVYa8H+IeF4MIpKe7AB
MaGmTj4Rl8xH63DQT6BjedYT1lzBR4zv72te8CaNoO8rGP4vj8aw6GjKtA/8TeL5DUBmiPUY43ZY
c6GXqguOGu2NQeMnAsmFJPJINi5AuRumDOVHGpuszNmyHrXL+oI3qfe92AnUVB43fg6uBFMtCvXN
6PFi6AdR8Qx0fa/jiRBYY09caqD5pL0guKlhEOjlQfZsmKpQABKuTrdrf6ln3EB+5plR/Oa05psf
19SwJ7maFTxHcpKRMv8zRLBOvQyBOmh0UmkVps3DJ5QhSx7wmDDyooa26asflEWFFiwYaW3/NQHW
hnoWJTKriGKy0GS1kD8Ys4fdPzaq3yVXcRJdUyslUN12DP+rjZoMlOOKhA80TpIABtcChkIkFImb
uLfQxmWqJdL7Yw75y5FLiFIaZYvk1xm5PT6N6gLzmXA/FGMIc4a5EqC/UfHOitQCVqZ0W2+6zhbN
p2qIylullGTNMMqxl2qF6qodv9D25PItukOGrxKq02cuyJvOVjnOwSd+1/SJbuYOk7lDepNXDyZO
exzvrxqkKrnhD/yVwGX0CQP3CD3VyNwoBMMo4KACp9oZelykL3fm3WNi5sP+3043fV9pX4tk7XHK
WBYSo4CFAgIoVM8O6FwadCGVCgYU1u0aTTcEAVPVqzUTHfl8y3ib2JJ5Nz/UmoPB4CHhR6ODuRjb
MkWA8+83TybWp4uPjUCEheRr+ug40hhGLtxy/7hPwoe6Fcg1zTWeecgLsdqpiiM740jJbQ9iOVRP
Vu0tJ1IhqxPgeTb1E+HwYvhlUBqcPCX+SxDbc/ubhKzyYlQHJITxXRgATTFSqAiKknA7g/d1r6mS
PPlyMobLDt4xBEfTq/cNtbbqQ5SYszl3hrJIcu+tvZ+8ygiLDWASLLjpLfOV3Jrb+Ts+8ci6iLdi
GFUcBmE8IGW6bkRICRLZTakb2/fuO7Dkl0VSacUE+5FS5kaZeJEMRtM4jD+SIuM9VQIvR73+2STC
thNzNiFxS/oFOr3V+bHm8RslWc/4nJjfPq1W9k25flTZfXOFovOzvG8GecRO/7ogPWrvb9WgZjs8
kmqP6xw4PL+NkQsbuVzkYzHSJK0LvnCw+SCevbMsRhb2dHeGtr0bJEcHOi9pCAfHbMVMSJQHIMfq
YsYxHPM4GTnI5CVArPIP6Apdc9lCcYungvPupgpLp04uyhIDUvxFxlv3A8BEWVYW0/hIL7iRrcWl
cR0flOikv2C4ycCADYtEwBT69SPNayPZ0QGTLwUEghMT4TDy5qfiFDOrmJB0JYPej8HQyb5zRzh9
HGjxeliYbZGpgZG8pWJ0v7wd+9ib51hiUJCbJF5sHgBOgVcwBSZaj4uHPFf8AoYPsSyVFCbHFgG3
i9Yi9ItN59ze6gaswalK+z99z7OmSwjXevBS1BLGs0EQp5ZmAGIB2CkInxR0CF22o4yiS9PGHdhN
AUTx5ogCJlEL0TXwGyF8zRBmtsr3AQ1BJMMhiXjGPzKiBiRGN4QNvMrswHpwZ0Dt94tJMKJYWvPe
KmgvHjMWrqOkCNgi3653N95aod5EDecqcJciP3Q7sgQrozLOH8D6ApYxpP+3VK21NKpqj4h1lb67
07E80Cht546KXUz+oyqrQjYgAeifqnwPke1R5wOjNL5KChj8QQEmHvsb3nU02QERQqVJp9MVTPqh
MhzzjlXQh6bkQvLPwofz2sOfJMbs91zLFClfa6aYUrRbhsUrCWF4/oarAupwdw35puuV0qXHXw6p
IMLHnYWT54p94TNRqU6Z4kISKirZCQQIm0J2rGvsBEPmZBtrLbshUcbft2v70mn6SO4QKUYi26wA
SRb7RsziXbcKYPvfkVFFIoSM+btsF/BmmmIAFYBRYEqa0YVr9B4YEU3atL+U1S+96X760i5Sf5mQ
bcZyP1+dlTwb7rIj6o9fKbtoj/zMl9K5BZ5dA7OCb3Cvj1pbL3sQnf5Tt9C0ZlnyKyWbF1AHEw+P
QbFu+R3/FHDEG4cU8J1kQMl6NBYXNqyp3QqbTGLnstxJXIL9rP8pdsKPfNL6vteCcOdu8hTxto3V
cIh6LTIcMqlR04T6cwBqL7XrFuI/2YBHPvD7iGLZ45UxKo6KWlhqI5p6s5HqIaSaYfX+N4kUJTDd
fGr6Yr5q2dZ9Im9ggN6Z2rq+nwFSeRJTDniKyEjsXgVcZAr65SvX1Xi44zRwPZHdhbK7MMx11csY
rRaiaCdQHBYJapB8pWmZqCl3IPv02TFxIE+ZHip0YeM1GTVOO0kzwQE7Irr66PVOL7y7/hLo/FCl
t10Of4QEQoPLbxZxn7PP79VEsRAdsk4Eu/s3HHvLpaucPMpgLb3/jFq3V77U74Fc18tdg9YBZtln
k6igTA4woCE5j0ieYNyhEdpEsBIRYy/GkUBGH+yNSKLRVlllJlcVXnUbaDKv31ThE1k1Z3OJo70E
qehzD4QKP3mfXaj9CAEHCIcWQFck5Z73mE3Ml3IdQ25uFB89V1Ao73i/RE5E5sBL0hLxMhdpQdBy
DSphJtFUz4LADLjHbdd5evmk5vxdDlKWboCTNNXIY5Ci2UIcUVCZkhkgpWsrsV9nOxwpQowgw8Rd
RrmANu3o4Xwmi585MUQ3kxGMyXuRjD/aGBhhdP+25AKXJq6EsU0NT2JrBG+8bDoYaF3b6xzypruc
vQbLrOZMq12Mqu64HKvPdq/8yscpwGlkCHt39NnEMAGG/Hb8TmlsBZJEhj67GFGkguQmswp0hNVi
NFbK2bjLjgUVk9BqkzAu7VyOZpxwleVowugqVO6QRBK4hpp8CUwrexAXHF/EEe1MV0jqJbKxH7EN
uTwVsBd6a9Y0QWngksYRY+KkjcaKvLESqwvACxMGQh/9y5PHv/kEqXtUHR4DwKyOkFWGqwtnxFzs
H9D4qcruuf3xof/5SBuYDYttxshqsH0OxsRR1CMCVE5eKanGoQlTpIhYhRbufjbXLIg9Chlj7DoD
kBJmHKvdQZ3goLhZg329fMyqwN6SptWdHofNwv6QdXNNaNjbCfGCRXA2RMI22tXfN9vg7hwPIN3Q
yzmKeUZKFW2KPY3TEYXaMgZkv/mUK25O0Jxx2hpYMxXGkVrhkP8Qbdv7LEsc5whRoeRkOLAu8nD9
mHgLRnmYMarvUV3p8At9zxfe/YsJxkMtZO1GjPwfYdPjFx/j9H+nm5iJ29hj/oBU74nbW5dIlYXZ
euspAVAkS9a6yBsxh+ncc+PXDZFMiPTkZn/TlZGWySCaGCfhXgdwFD9TBXk/hkEq8Elvzfhk3kMV
6H7iLDWF4QBHhoQLb8pmj8nWkEpJsF5yQj/h9Lg1VImiL8R8uHztEs2OQco+Tn0+or0NkJ3zgtLE
DHyQQj6FLG+wmpO2RrWTjnMUAjNnl3rfTUszsKFHiS0VmxTYa2t0GvVfnCeZIeJ4JDQ/BtEOA/tT
l0qYvPEl2Uhk0NRMhWjhDORZEvdtJMc8rCqeWoXBbfTBPBHQ6XtMhPGjMgjzmoLYWPU2WDAWwCd4
pCnKKDH6F1uzgyWATh4ml/BK5xn5pJTOh6zdvTB2KUAA3PVU0pa06kTIv8xboYTdj6iNidoe1/Xj
UM4KKKts1lLGoZRGS/rlJsmAO8zW6cG+xAGDQo6stbimPSuhNmyVPfdDSvWjBPDI1TDAobSuUqzz
0uPqYNrDnj8OPvA3FqAL9X6M5fJnCySK8pghE4HiCk2lu1mvo48a0V5x01rN5WW9GvO6JYAp3/cw
+NV681nWCzPWhAcJa1ITRYWWPO/+Q8BLIa+y3m4nJGE7T1y9s8RuB4vweeQgze+FPwZCR6rL36J9
jfJSBQUEbtoZyfuLMxs9uCMoKzmg/TSxUiqzY6qUsoXGrL82p4ods46LPNQ4uDLybNQhJ/i73h5X
8PE1Qzss8bO6JVb4ErDntur0lUI/jAUJchkVhtf4MWM/hb6X2dikAXErPTiPTQ92qd38fyK85Kkl
j+eE7d29zZ50sydeG2URy9LfEamictXn6f+1/2dtzx3f+eiF4G84xL7i1kjQ7778Q8jX75m60zk9
UP+4//U4RUapQWEKdmK9SYusfcTi7G8D5mZNrtz+bFLbUInEvLJo3qrwtD/IAsCCQuNQjo5/vff8
p9xt5m14Mv1JOF/1GfT0/xfiTZ7XQKi3xoMJ4XpXN8rpLNpPVxHBCCIcN8Vd+ysHo0m2/2jtMAyX
TduLeuWGFHs0ig5I0u1XhgFKQfGSSHGqXSBzg5gFMX1b62ZX4tHYTM/rXrze4a6MT0Si2c2Mj1+D
Sh4Igl/To+9qIiG6LpxRw8DB9HbEUFUA6myJRWreVOzeiwsY5u4IjkHi0xFCXLER6/sU1pMKiN1Q
lcpaNb0mW2dNGmjjUtsT1ydDw628R1lBjvl473LIQW9AI17s3tf1PqDqWlCmSPHfGsWhaRhWq+gp
bXMAaj22Qoult3YdQWAfQ91jweJzvY81MYbM2a2UbMWriZ0MmpX0vYSlD/SO9O0vORkaFalGH7r8
y2Y/tquHMNtkq3rCK+K6nRWoUYwPa2vAmpHyNDMMnhQrEupoRkcyp7O9XjyWbl1qJ58hhnTs7R8d
lqGW/erv6B7UWvSzd/cIO9tFVFgX5nvXZY3oFf5JlJldCmX5yjPxqIBo1OUzH9fELH8d2P2xvJ48
fuqGzOfQT5aYHWXmEKbrriXrBbmxNchp0D4w/AjJrYXQKlfhliwfUtGzNAciC2Coupuhg2TSKAk8
BXZz1Hr9T6rvP16Tx8NN1YIhrSAbql+9goyVVQq1r1UTnv95e2rNF0Ca2sH8Z7L+qfk+R9FVeeiR
qM33l7vRkOyYe9+nw4Sj+XYfGn/r28byBxTT+ZrVxiFHYqiZ4dONnDT71t/ecQuYKqJz7bFMWFRo
ws3nTxnfi1gnpm66V3f72FbxtJZYWUdDDl6clnTZpPjPOwFu3gukcr/eUK43Vtm5tN6t82QqyVRb
5eo/XBDUOt2tgL2laE+eB7t/WjDP4jirHh4jnmCS3iG0SVbHkR75smc+WbblnupX4qO9Cg/l9j0j
Cl3tp+2BEkC4qN+0/Qwom9gK3VF6aYrT6o456bArGDgSax8Yn5zjUi9NUoRRodsID0SWJbB85kph
wAc+n1xhnzO90mESO07ZpIf6v7YevGUuy8l+5z/j3PCHyinoT5XXKj+bRQ6NpCJO1sUjuQiuSi/6
eRBLpCdL2/71FE0VWSr4376beta9/Q3lJjbvlYSSooIMbLFiRfI4M93PD8K16GIvOqBRU3WrBxGV
3Y/1rl/XByyLGcFqtHrDtKyxxLsBjIS7kCpV9qCr7uGxfLwvES2QD/JuEjoIfB8aKEUSLh2c6te8
oPWyPHG/PYJCvgsFcjOrpPTWa0Xh3dc2xoAQcaquy05UJq5eXYfXm5n5clc4dtYuOE1Elm1j4ZEv
U/4iSd/2qz//AHHSNlxlab34SSLa+E2eLAA+/nBDULOjSP4l1+7r96SBFcW1J+KcX6+5fCVaQEqa
ftaxrM8BdzEsuPst9cG5KNitMAX1e9vqXHznz0aQwxTfWhp1aK0QO6Mmi63NhY7WpfwZE6m+UKVl
EaNiobgrVJzibesm++pEyundeUwymnzhEjPphs01BuX7wXzUq8hOYHOpmFJ6AajUN9aUGyiKaC+4
YmG51Xkoc/xxtu4GqKl5l1BeJhJWNbeKfhjUbvYkxxPc7JFdDt18vAIWbvT/f7vuvQYQKagf4OUG
XS1AGtZf7ieo+lDx+Es8qDMwduJHPMjUOZ6w4IiAL8Xk9MYTJw3PSD3+g8VCp3WQcSpDABByZFOo
sQeqAWKlOH7Hu6V08PqfFzYCP0r3fbrw+PuKPd0gNZk/d4Vt8wcb5gC20yPQvtbIruzF90cl6qEj
XJrIquS4qSxVtbZ4h14J6hljnULyFtjrgU86mIQEwCHC5xhB/EshORo1Yh1nz4xLXfG0KY3niCNA
Kf+E7jdNqgy3Ew7AzVd10pedlvcV5snUAO+13X+UPR8gpXkfbypJPKJUkphT/6c7QhhjHZcEC/6n
/bWKHxCVjqSCfWeJXnOv7groAMlg7JnoLTHkkn3lci3OvGXrdlcmX7DuE/drfAdPhF16gjbpYbGf
632hLT6UGda2KcO6kU9jhkEVfzXTx68Oiscf/GiqcHTu62BOy/4DgdrzyxMIvXApEu5LO8fZ4YOn
hy15txfaXZMqB8oFQnOF4Er9MiuXXX7s0Q2fGx/NNd1RMtVq7b1oZX9EEo7+Ys3wci4qkcFnCBTx
BMNyA+MUyRIH3PGHoteLcmebeinit/GpVCCf8IZNX11E1XchdR98tuYTmfsH6ClGpijIpJXd/QCP
RAvctbYGhMdOyZs9VjuHGjZk4sJ/knDEYamz4mKA07BP+Jt+Ol/587qxaP1QalvceHdnCjsSY8u7
4gess0zmqO2WMcITiGRsH0XuljWLK+rIbhIjOJuIknfBEJ6fo6GxBxOB41lHuHuq6RS9ibOdOSw2
FwQCTwb5TeRs3sXCiHcIpo9eHy6XmOKGV8SY65HSU4q7sGfzeUcSPhqmOaCoNa4Q4x48Ac04a9OL
6VU7oTiL1DHu3weAG6TnlnVWIiZquUizUSTC1VZNNDu1NPU72I0lWZ1Qyf4WdRv43LA37o6ZngfP
ZVFSTdKWjXkThkhryzvRIZjn9l3O9h97e/5TQ1iuAuxJSEms+8Nyad6hRGrUxZmK7zBIjCpoZRf1
wJg9uCtJpUwgOHfF0DUDZeM7NJAF2dOn6HmkU1YC76k0ITFyaoQIS0ZBbONqpJGPDlqg5wRJNtGe
a0Brv2y9yp18JFZChmCiYXNNmJsEyEOI7la/wExQTmYJjz04XeBw14Oki+jxhfqcyCI4WJuK65UN
NRM2L7FsZ+Fj1FYJRbjMD3T+jIrhKuj24KSzpuTi37GeeeTsE6QiVfcZNWuNy0DGFeZgIOivAeku
ZBk1J+4elSzLWy22PnukiqmtCUFxOIBuATFDca7lQbctMYRFzFMnfzdkD7liEEoSCDVu1TJWaLVo
AMBrMiDD2YoFnFgnAQkkyA/tdeQ/wG2C4l4FBmRuLndtQdmpaY3ip1I/qCbnraUwVOHCupCRKTvS
ZUdxpY7jT08+6yyP/+fR8d+hk7weqDo+COxUuZTXtaeAjIuEfYcKydu2GzZx/DloF5qMSCiVMP8k
vgzCIO3GGx1dmmn6wzAbGw5pIZcJwK25Pge6Vf4UrBrwU4BEcFjB4+pXHIT5Gl9n5G3+eMCX61gK
12dBfd6+RdZ2KvX+emE8BGwx5ylVYVA5FGKlfGb7jVpbpAl25S+ooP53cj+DyjMhJUO8wVne3cV9
2C0fXFLG8pDZz0sJ25PI3Y4DcmFUWo8f7psTrO1Wky5/0qMK9U7hEkEhzQpzcQT+1ZKKssxQzEN+
uampPKaQqbaJwS5BGAb6RRvXSkgtphuYPnV+0lxwAsmgDevUC06JBdb1w1aLCP2ffz5IddyD4f7x
m5KdU2XGLyf+yAH1RKBAg2sQ+aKmkBbAEB0pUICRw+KYypoT5fcbHqnR8t5MpuoxgsN+XxEkF9Vl
cKG87LK79LQRmRPqeihSDc8DOne3GsTnYgzVSJ/SoDHQ9IQ9Og/brTBhWtvJcziUwsABHFwjQjEp
nnR1C4qnaPLdNIQGtQ5KJtWahHBF+5s/nDo5Cf4BUQ2OLfYCxgtBzQtGJMFvTTEQ+qT0m32QXo6H
MTp+PVaJh0vUSvggU3N2kN4bKyu/MpGsUg9d6k6h8Re0RTagaUwBENDblLQcSDlNTmcJGRfxxjf1
jH7n4vqQCaF4v+hu46N2WCvjhok8UIVqESWz8TjVLkwGT+qHTgAfDAzMAlNlMI0ZTaHr1GRPzh7m
w/f5dRJkG5NnyWU8NUHJdrFxVsZICexyeoyubAbxo/1SUHA1JaWtsqCPL/lGjGoBMAFTUnyaqw+2
rSYAb1bgC4BnMKyx6knAlQzzAZhihnnaFH9HaAores/CoDD8dRgWb/M0xv4Ih15S2i2/uXFjZLOb
JpoEet7P4CrOjYvTFupnh4i7YxskvgarbXGWy1epvaxMETMQxcUoRyZxGpD/eG+9eJy6y3i0Uegz
2/G6FMVqYGgm2L7BiKLBmC8sVbZgHkZdXsEonbPaVWa6iOliGA3nWernNR2WdzjIkOec2nDpbKWA
rJ0gaIY+q0ISTAFHrUkrjXYEEEo8K/prGrYHHdFDhegeEEhSs4jFVdRSWnjrPJ/GvT0bFmssorPz
nQW3MkXGr9GIKzu8JJZSxAalnGi9t72t5ZhqfgfoDAU0CECpUWaiJIUh36R9HvKeAbeEQnn0ucNd
VoeBELvFcCDdI8n5D4It1HCU8U3edXoVAhmMNMjhbd8jzv36CyrMe74cnEY/kD6huwTr98XK92ut
UHunKuehRggK85vK7avkAXjcoMalEw8Xj/SG245k5EUjKRF+Qi9GShyUdAVEhXd8YyZiFuN8KMKl
XKVojGH/XDCej2XNv5YoW5JiGEn2Uw5merSCs6t6BqnDa5Aui5Jw0FvISIeOeVZc/Kfuls1NiS5o
RZMAs9k4JUEZQnez6VxQqbiCzeXjDqdQVD9HsoW8CJy8C5B2ayLVamsDu/NuzcV/Q9bccMj0uELq
oujr0EkiOaijp2Eb2PvQ3wzRT49oTTsS4x6WsqpBaXOYFnYEQW5ooKnk01N9hGbIBT9J20oBHH/B
+UO0bwSHLCSzYGRGWS5i7zOUMG4TQKDq830f1f1ZRIsAt7nl/YZMmuLNnzTRCygIQX0LeWpPewez
WF2z3Xe4/uV5MH+QUB1YMyzv0Rq/1XdCCETQlWQXVAleWZXzOhyru3XgJvkeNN55REI7+8XrK/+H
NmJeaYnu8GMh8pUccnPkzj4hNEPavh0VzJoUZUr9us9LQudQkQ1QlyA9jFTetKuIS8A5+VG0MvEJ
jN9cPBUL5f459YkTkIxJZW/X+PrS/N1IhaHPGxXUcTHonqhX0HNB9kVINQJIVj0acTwRTWQX0e4N
NYkM+xkpTxd2xq6OfuFXUQxv50KGOyUpnBpfzb8E/n9pI+5pE1DqU3L78sI4zaz2AMdOKRsZYhci
ltttXxwAO7Qn1RpO/LH67KDo/EHw3WXG84h6ag2EqIgL55qMeO4tBy+2zcwoz7QHgXmm+0DUM5oe
XqDkVtBXwQqxChxYYjOez0RArRwbrjmv3xAhEr0m7doMThZBFCdJ2A0CGt4CsJYgoBipjr5HJ6It
NX1vuYS6HcMxpZ4EkdhpbPG2MiueK5LO1znJHZNfarLTvFu7ZgOVMZIUj11ANeefR7kPoyGSx5d6
+nE0GjNLFYEDx1tRRIUCJctQAy9wwJunc/biMtAs1YRKCrJBBvutTQU7ZCv8XSSMxwACdM9aFaV4
1Yol5h5JvcJjGMXEDCrcGuGgwJTszAI6fonqrHahz0t1VSBmh6OEYKfbss4zMJ3xL7c7S0ZBFfW7
E8M8iJfpdR0Xy4mqoN0ta6qH1+wMlsMANpgWe45Rs5Pkr2TYDgcMckggATuXs+dx8kS+wMArQUc4
mvT4/LhK0c0LDtutcVqy991gc3LLsholXQ3kLd/t78Fz5sKwpeitfix/+ltCc2hQYoVw2qdwxHdt
FeSwiWLKaPGt6tk3B0eNWJkb2pO/enRLvFFR51awfAyF1yFothPdaMQlSZF5HZLg9eFQMHRZWgJM
5RI9pCDbGTY01W/6xQE3ycsST6SlXQXAZwUxW8NcHpAomN2YHPiBp3q0FHizIgmy0KB4cTbR1++h
ZOtjFjO0EC0OwZIsZUTHvMQqCJIvhDVowFABlfm4DM/x+Ztoy7jpS/Ha4NDoSa51PdDuIc4sa0/u
UHKGBKXjRpdC1kQvHznvyUFy0aUIXtm/yd6cuf74QPdILK/qJEeyFb2pNodSsdoF0ZlJrFCo7rNj
DvW1t1kmm4tYCVF4Pl7AUwqNc8Jq6ODHbuzBIqoyP+Mkgvh2LBJMY37ZDur8qWbANl3qnOhewNGq
pGdjUa7o3A3fmx80jVZQkOBBQKHA1ts5L7T0Vy6W1J0ZdaDdChNWfwEjJRxSbT/sNriKfN3wnblB
5jIds6IKQ29mDiZbrOTt70RPi5Zxd4iS/0Fch5qSBO/cSGy3C9W39+ubExXRbxitZPkGF6y+s9hP
6j8LIwRoIPBEYMu7FEGZqJa2dRnSNSd7i8UHxQxcdPr6VU809YZknKLVlOyqBsXvD2MHc5WBj8Ic
X3McvdOS9YhfB9G6Fvob4PsuZfw15Zo0Q0pImZvmgM5ssEoFe68ZPkOTNHRvxx+jGriU724CKlqC
b+rXws9zsdW64aAzRCzU3k0K83l37nb2yJjw0bJt068r8B58u2+69XFoIlfUUNSw95dE6rCoYFe4
NF/HNVHIle9Nh08+pVL2W8MM7SU7N+IE1wqGvKF8AVkMi+/n2l3xv2s2krdswaiT+rJsl7MeT4Ro
cl41eR3JUkJHrxO6o9sc0kex0seUNhG6ZQdAHfTaL0aY8DCj9r2PVGAU2lb5GFFc8nr+Pp47Yn+z
9mYsolu2tSOnXEuavuRdy6TkjCfYUjLsAoom8EfJJVRTsBETar24UVzLubaraCgTxDJNxST0pC/I
v9+dxVv7VgSz9Z3qrf2/78BU3+OmvUMFcPqIZMlZIkKp5ldUMZuEOIO/beHAJZVJpLAzbSToy3J4
Z986PMeIbXpWYhIRLCulzLEzlnvb55IsQohMxM6VMMQbnK4UXw6x/UYv/aATAsgxx27U2N2hzNKn
U9Q2k0+ic48TfJagA+GBrwzDtj/dxXHosRgFAAZLzKqw6kpA1D3cYYFwhLI8oiykWci0wsyq1uR8
cgob1Erjt/lXYP6PTdwqBKKsDkYrXYdhy5K3RxswAr+O74L4W6KexMra+UpPHkcc4f57qTSNKVcU
3ccSuQzLSbXfG5mJYOLUHqvzxR+tenrMybzbc/daCqbP1LsxG00GOBznlnJVL2sni3edPpU4yt8A
+llFqdCkP8xIxr9BxqyOBFuvNrJwJsUoxsPtitGoyPKLg6QFyRoNdbgRfFALPfYu7NxlWeAMjqVQ
kc5MB+5/in8EzFPL4C/BNBnIEZvBadUhLrhPxbn8jXoGxn27j3E4S/IVASDlb7TyBmEyltFqXyP5
/TzDfkeP3LOGB8O2Fr08AW23yGh+Xe6faQoj2hplNWhBlKW0C9ar/IDnLsmElEYhvFCBUPo/xVKe
BPl2Ku3PnkBBAmjbkoLgSus2fFiJURVFXTc8CF/x/lG1AXcEzmyKS1zgs8yMOOb2u6/z19aSaXEB
Ui6PPfhngtD7RZyVGrngoDXe1ytKojsnLNiVtHU5JKXPRbEXAiXfQzmzjoYYbzQ9bKrTCXLYme8B
G5Nw92RUGcy87y9jcEwOWSzQTsIQu9KDm2im68rmr+DuZpCQDAOCkDO5z+ZfLAsbRh5jxGJohDfE
rENj0EbPA56McE5KTpq1XM9VhLryReKLyicTahGA1ls/waOgzgI6BxFn/ftUOt+Eb6G91ovZrc7A
OBVz4v+kiPNx7xURZNCMIiZZpSIqKdfAqAuvOUXv1M8YnnSAvacJVHqAo2NuJEhch8fAsOcMXmFj
yugTmDxL+i9dMoLtccpFnngiZLDZHURAQVq49pWhe/jpQAP+0CKe2SdlvyW8tM8uWBrHapnJGfEq
NHuDZsJOcn1nfVElYwZGN3ipOCtpMgi1b+d1Oe9R8KBoxT4ROiELVnEP9LOEcLnq6WNP+jTgic21
48gA0+QE8JrtVxxm4kinbano/isNkyaz5xubD4vXXF79gZmdQaAwzmy55cSGBzxFB7vcvfYpSvfm
ZjYfTEWBABaDEqzIDEYgcCss7f0lRqNOUBAt2/+c+uWG3PbXilcosOfL+ibRRdbY69CTKhX75lm1
sQ4X/blGxCA4QAMaalsoaIUiylNTta/CUSm9tFEOI/FBSvgL9gSPJZ2Jxe4QcChL2V2E9PkRpVrA
RMFKCU09fOsDIw5TJ7VnQYcoY0V/6WENOeC694qm2MuAY0qU31DxdrNZcDoulOQQLiVag/h+kibO
YpESEcEIPqqcED4DWsoFypZDQBVEw8Y0cb3OEfBgtoSlVZxz4BK+DN1DaruwePHnZ0Lg8MQHfSsD
FemYmZGXyURp+AFvD5tTYmPY7ZJd/of8sJ5CZ7f60l7xhHIgxU87Hw8/OlUlxpOmlduJvqacnH9A
d536LRqk7F8rqShXVRhPGfuu5ZsxSsZQIGlcASlYnrhnP+lZwlHyaclsi+frgW5oL0XV1nd9+Yg5
NgDnqPNTuKW84pRvD2vsHyiA8plL03mqAQcFw5khpQPoSDT4FqcM34DOS2aW6Pq8P2xgPosWYoOD
ZF3zm+a3Ac1lBaVskohuz51iDePxaFpmyv+fIMcAIzjcB6e55Xx3VX9ITeVYI8G6XvB06p2eHEXT
0gDPusY0C5MEMN0xAoLrjE4i4VlQBP5mh6JcxXlZuOb5/21RmNUoN23hvUNRFLu2RribJQ8izPWr
+9vWjmzHa+8/MUoEUutmDYg4qKQQGthLBi1RUOT87e7RcxmAZ+Ra7wVU8QaCFw2+jxOGm9+Z6Zvi
Qf/AKefiHmXGaoaD1WdPdHNDi/ncFP7Pm3Vyj+sXRLQD1j5AYMrTQA1uUY+HRuNYyFENSmcUlomo
otyPrae7UlCykXjPaC6UeFWbKmjZ/4005rP1hChQSvn8vPSQcRkaZn2avMHSSSI79lRo3/6EOekO
blH++8b+4zfOHlzvUmc3Hb2n/TaVTfEqI7/T28a5avnfsZzkBznCTSohLCoAD9LSJOxLTyr3mZKt
tWbdVflgNeW4JNYUoqa3sB0d3NVZYoQlL1M+tLHgt4f08eC51ITuFsqCh6vK6S6cmH1fc42MuzeW
YphyjHP4n7TVsTJjGVAmuFK5W7Ygeze/kVPu4onxxxYpS1UKfOZamaT+hQlO4zJDXjcPTF5E+d4N
gzfdQrfV63qFhPDFT5IDm2W9UHo2KNVfdveRS12kJ8Q4MA0rcy0UHY2uOceVplELFKusy6+pDyQX
N2L+9PlfrQiml/x5JnLeihehnFJheORQNGfj1uYBDV1gDUqWiX8EOoLHBvimqYoHFTL0wBBHFbuO
ZUDTCM2qpdFusjyOqr7zLb9n6N1UXJ3uKnP19qhTQLlfIrbfLbUCCJXQP1qIAIJ+9O7z4aGJ+W4m
lmoFmwxXWa/Ezd0yQki2FMMcX/DvxWtSAWi+BAnttlh3fyk2WCUepXviNVePYVdydOLFKLYiKs5e
UoyR+faTkQ8yk/eecB0ETK07HeVRQqVSfc9hmFqJDAdtH/R1KHQ5DTwSL7dLBtiMM69YmAZ8JLJD
/KoxfIb1D/dD9ZN+ZJP2P8eX1G1Y7+KIY57MzXddoRZ02PzDOrHWpxGDP1qFznepVXhzlqzgESTe
XBwTHoEkIV5CZY0ymgocxv/bwDO208daovG1AoDdSpj2CG/RbUqfBiM5FOAegdPZGhFeZ+GOXyX7
YRr5Ou6VLPIUmnk6GgzcutOLXSP2NoSmcRFtYSsnrLAHimbnhiCtBKIAIWrXojoqmvMB9NhSSmTt
xIdn84O1Oo3bxSXEu56O+iNupvwtAyY5MPoyl0p/37nHoolbppEuDEm6OQ40T9fNe1U4CFXEJnDw
EpjRvNhkkbTkzW3/boBAir1P7wHA20EUePV7dshutmAfYvjUoe+iBlCNd9XuNqbeS55nK5JXj6Z8
0nclb0Aa+iZiCDDjvj+3rc6UhDr4NcLZ7g4v0G3XZvuVIXRIfPXkpE5dhvj0tVK1l0jFxJM5jVEK
CgTgQsgj/rBOuZ/ImqNjZA+HjYo7a9capLlrQrDk6yDOApBvNrPSKopxIVJrGV7xMpo/BNL9C23/
gaMexraST19TpFS902h2lLYA/gHDVSgQYIVl4aPtiOAHhcU8VG2WBDzn9QeNL9XvNQbbr7iF02Vo
f4nHD+p5riU1AI1F/1NypUWrl6ayVLPmaeNDF4t6jB2jxNsVYY40XRd6tjgzb9Z7Jz4QUPHxoJ6Q
XCtYb/A1aKTa0fZxZ4xjuO8cF7sSZ03IIPREeJf0CfD+kToPUWTzipgo8Nn9vs0I+hRlYPrjvhdi
xi8fc06w1cbIlfhR9bSTPyc3s9SYQbfQxmvtb8yVeP6H3tVPkWvauG+pRNdH20I1U15TrAQNR+74
5ZZyBTgeDnCZ1hPFoSe/dq5YJDO/JfaEMMOy1LAdfzUXn21B3rfNRQB/e+gmQc4Hy0Q8wqFJELt7
vaPceUxQOfe27tvoDsErGlBjT60x0xf0mAYKfEtUBgaZglkta9/oOCAryTFsXeQoQSe8X3fZYuJd
qUhxxsv/fXzNZFxkeU8ViGPy+zuCS0dRl+Ycu00OVXVfoljRlpsfobEQUnSER+eSjalP1tZKtD0D
SkJFrZK9Ku9DXg1taGeJ6DodSGuIDNhkjCwXFNpjklEPjNRMV5Db1E2esUnoj16i/ckdbtOzaExh
lZYzD/Lp1GoYocttfwnxqQOzjt7fJNthLFOeo5vcrNxfg4GoW3Vo4umQ1lBcJdrRLIORPhPOgYoj
u33/1s2IDoUuMqHeJ1Fi9PuezXRrvdEhkgzHpZapMlcfwq18C3M26NE0T+dAK9OKFHWxcST7pME/
zguJNMJmIsOtGm1LJT6rhyn2jGSjjCKcIX+HgoiywaBk1avV0erY6OV3TSNL7ZrlWUM+hB0I+Bzp
CwxgpsTIDBN9sxqGy77UVEnOERVgTaODj+NeiXdighEwKkfmCDnRSByjhRsY78Qvfp6ITR1LT2KG
o+1tVODKwLoI07WRBo/IXUIW9grPKWCmD75uWt92H8ucjBvEBJQEsN8me9vU+1K1Cn8uzlFU8e5P
4GXsO2aP+AunPAhoinEgjhSD9db0slY1DqXyfYOdjyfa2/TRr6H8s0AHmmtqqmcU+c0G1eqLoxs2
ZgSliUH53/i7sbf3Wx5A18fSXMxHxsByzkJ9sYhLTFFUbAQ5V5NmXff8t5f2kqa5bxVTLMRhTEHb
ymeq25N7CinZXeH1rgdGHCL4oltslF5g0T70f/lexuGfQWzMYij2B9scrswGkNxNKbkbHGTkGZTI
pEf2TBSsaiH/A5xCBdifiakliJ8YyhkMDZyVgYoKcs7o4/AZz+jOj8xyigWGxwT7PjIEqo5pAldv
RRMkpGBo4hC3J2zMUiS0zqwXICZO0jJZpqsxxG8m7mFvAk0UKrjEDcvIE+NnJf9nhTuRAenu5kmC
NEqkpwwPmTkhC27btpgrgi5eXC4kIMQ0PpfFijpD5q/+27jJMZiupPMFO2SVmTPzQcLrgx/Mi6ux
zyELh+X3Kao2IpIcn4EEiPRWAb0+YIyZxiFBtWvsDrb5BxdE1YCkb5fYziuqsihaPw0adsDsM55T
j9BGTPKlgJkoYof22wdR1Xq6e/VAFm+9z5va9JM8clkHIm99KClGA7axV09HWspPS4KDXvygrChO
78GVSIDEAtq0DpwKGlYAwJbDKluCjdM+8B8sGsBHPB6EFFynOeT8lMw556nTyiBQBfAn8Q3GEgHO
UEKV80BG8P2ulZwKX4R3cFpEUtGADDJfnbGjY/eYAQGvE4prkQSNRMUwsU/JKCeNjnL+/zFzYucC
XxvgTDkPPZjknEefK6D/Qj+VAkZ/sCJNkjSAjrVhYHzzCnyfxJ5NJlltsqE+Yh09Rinlxe1jmEVD
viOXFWBI5aiLXfXn3/Jd0L7bGeEVLjBV4X3koZ0IzyappMROrsI9sfEnTlA2qtYGiilYHSJfinna
h2rK3wHiD0Ow2g4SOj1h5hSRZtgJhQBxTTrOew3pYYBpbzAsDWOy4UvIHvl2DlY/9tvw+291Mzm7
ZaJbtUV0LeThjJQ4nf+7Ytc+burBC9l97jVCmPVYsSp6UtN8QcCOxuaH9gprRvxw2noSeMhi8uvY
8WRklVngjKwP8yabBE0F6MuaApMb3f1FgUTqdpweU+2j/mcnJUaGj1DD4oHij5yzMekFEjCPElLY
C/DSyHhg0s7faPgQYuL7IB48xO7EFzKHbID9x60bXlI0EHaWlXku9EI40dVlDzqXQz9EAKS8jvNN
qwYZIeJ2cjUwqHeEDS6+KTU4H+22NMo2tal2Zgx1zKk1gj9tV3slIs+LTLyn6jqFRGH5Sd6JuX5m
ICpQRWI1GXwLuMvAt7Ke9grGL/m0zYnDvqW3lCDQOL95tj8l7uLgTHE+/6/4c7cF86U9GzRXU2nZ
BAmfOAM3T83IjAm/wbumt8pT/PYRF+J9mbHa4KvCLURGC3vQp9cQ76B/3GohOB3eUd8B5ZZWhN16
IkSGvujSrEjnz7Uk77BCj1eZxgymK6n0wGm2G19Bgdz6OMyui43Py9G6GouiZAU0jKLRbov2R4lb
54d+FbAS7jqQFf+wFqn0MvgQD9QAuaGCeFf7Ay0a66ea0J56D9EnS9L4rvKrtdLQwgpiX/BELkiU
L8EcA/ZhKHPLMQni5HxV1Ysap28gY2ITymOFWy/YZ2sFvnXgZJDy+qd8GaDJ25SoUYSB5vqGyA09
H36xY4eijmgFMZZ5FCQJBGjUN2+bs/mENGk6xtg7qbpVsMaZDOpAkTD9BpT1FHI4rUg9a45rVeZh
x38eZ4US4KbXnMFVQQNgem+ZSx4oNQR2bmQ+1CJc5P98Td1Pka/o//hpkB6SFu8+sPDTRg2tT6bt
GzMUSIIeXb8iNiLLBJq4pqinI7Vghg9Hadan+kKdnmk5tbrvqmHkGAmzdsZ+shkMAgLovtPnwYdE
Rq7kfu/aDL4ZbHh2iulwRSjlDUMdN6M0sRnLqiJSdPOjT+y6TR1adLZDfKIMIlrTp6upTnibzloZ
YjLDz6v6y1B5KuMnfnqlVF1Rf/U7O1N1C+aSc/petlzL3fyeDCVBDlDFYbjwOSm6PU35W070T1i0
6o3ZW0gWNsUklzlCwmUVHrJVDdzRuw1Pl5YZ4FXkni66G6To8thRwvauabqzLauRYSpG4vy2SJf6
BMt9GrST1gL5D0cJrhFepKVmLVnZ/vFO91w7nLyOhLRr9JBU09mnqS3o4c2In9wMYtS5vOu3Hppz
3nSNi+dId8kMlpmjn+FciN6zLgetcZIS7jjcz5IzXKe140EamwBuBjYFcuNlqXSpIzvG3sYqmE0z
8MeRyWYaF9CJJfUGDEcPqCGimScBxgarL05RgI4KnFreOOTApbVUeiaRp6sodUnGxZcUpLot8W2m
8svx/nRcP+UeP0xWI4Hp5iKtmHMtWg8J1NJMB+D/p9jdc940HfdexLwlaMPYcf0LT/tqvEw9W1WO
9qODdr/hJXgaP2LqLYA4CVrkWcJVtOgpE62QvMs5U7z+WKAk5UINGgMApmiklURK5qECky9lHDGC
P6v8oKub0J8JMhcFFjR54C3WaIkWa29SrQ6s5+1AM76J01F9jC98X5EqajXUVVSKjoGTlUggvLRS
2med1PDQlzJm/rRqIDjz33qGGDoPuzmmH3MDWLQGnsBSuAjL8rsLSl8+UA6+xfN5Ktn4Nby6GvII
U7kd4RQ+lXS6qHS+qe2RZFDDNSXxVnx5o2we3uhFPmbI2VuwPkfY9UUEqVdRzBUXrLTZI70znHW1
Oxt6QjOERXutMuLyasseT49vwLOgoWQ3jmrHt98S4bcbSlMIBfYpll7ZBJmG2yyj2Tn6al0hNeDD
AZIpVRTNa4m+wUomBHrRclG+cHC+viNUkZazJlOt+/EcEn9c9TFGAKAaXgCQKIKQe+qHJuDBILuc
lnDrzg+AfMcU23rvMs63g+A5TV5zzGcARz0edGWcTNuqSD8wHHNRXuWfSzp+OpXQ3zy47W6eqP/T
s9X6gAlLGH+4TyESh481o1PhoRkPYr8Md3AuCnY0qfY/nzL6UPi6U/ECkLj4jowk2F4cMMg6627y
gD3nRGsM5CioesSiwfyYFKUBz+3H5gzlbKUMTseNqZcKHgKxD6rjsi26pRVR/rOKnso+sH6YM3Ax
zrzp6rVK8NM8A5p+zoqUgQoGy/pu/GdQaVohOTeyVz1smdafEgR0LzifbXMQkXAW1pZH4n55ysDc
yjKKQuzC05p4Ra9066IkyhYV98lvo+DAt32VIIe+XgmnbT5/5HkYgbAoynwQDzaJY8BFhu2UaEr0
IPBcbiq0moPQGH1pJEPoIL4yAcu8OCs1LXY+32nPhPj4W/BofPTxG/0/JkepxVo5TvNWW286jQuJ
mFaXodge6/UcAnoAJX3AsNj47dcWmppfwZB/rkDdlZY/QY6jCu69DTy9CvEWcNsQisvsDRrZi0L+
ueGX+UmJOsi6x4/DuXzWCXjaXGE1EXdIOO9NGvOyhVLGkdBefrA+SNm3wrQPf8YpIqVgfUXz1zEq
BQ9KiXmhqLvVtcM6ndZv1ujSVhrHFOHUHpsw2dZK5siodAoOiTVx43hJvgrN2nUmm9X1mvAB6gJt
He74SkuJePbj3HT4C77nU7cqFvmeEbbmdhRFkb22/y1H/S8Yv1x5RycIt5AXpq+zMb4jCeNoe8eR
cQ4QKmOJWqOlrjgSqYf2j/AAaU81FpmKiHDJHKzjp65hkI4JNLYY9Cqi85F2HZGVXAxQv8V/XG84
oZA862KDAkL9PNGnIQhI8YWQy8O9pzNtFqCa0NyJQzAvqClR7bAWXs+rJNLX5xndzZYOq3BOlftQ
jEcZqyPUQGWgtp+eGurWqX1tAsWyZttLI3JkEuy7U5+kcv0v0P0bWnkYbh3kLP78ytji6DdTrf8L
HiK/xQIvOqMfhvnB05ul6CcbEIUfl8XuI7y8pVkzBCtC9l0Hcy+PNKEYXO/k+97l4OGOn0A9Nyff
rf9XwIlg+zLG5XSf7TmB4mWXFWYaoC4aYKpyhq4hWfVPkQfZE0IfVqxDTf2xTUBncL3fKFw1NcA9
WcYF7K2bDMaWPMnKfFg/7D/tKmr+3dAILw9CLa1NUAKKXDWa45ZS8Oy1ixCkQx15rhTdSnbpnaSl
kmU31obxmSWr6phsl5C3ZaLIwqueYc2K3tFLzPel7WCmF0qhTvFW8pamXLWQeM8wt8ow37dDSh+w
Ka77L0G8SEcTL0rM1hGtg9Y3X+L8E5azIqJjWxAoi6oxl77D1m1Wdc23DcKBhOVzuk62J5iTGooS
HSXLsdj2u3iEjZ38bVgNGRQIPY8yAf+qPyckCFGqTrMRdVnVif+SiiMHcqNsdO59urd29AHCG6CQ
/uyS1430bG5idI+BofB5MvQrfJmMnjjq9mRISJELw4eTfldlSKd5WucTfcBS5Is1LTt2hSGnojg9
yT263F4JnyY8mCDoUWM59wPbfqwcPUWMK3TeaEFP+gyS7ajZm8/nN5HSW3NEN3t8hutD9CxYAl5V
aEVuEcTKjDo8jlla+0GhX+4mSxZghxnd+uA729TJWGiflW0NYSx4kwHC83E1hwHaXTyms7eP0LuJ
FIZE3gXtEIYgJf9tLg86ttZ6k21Fgt/iX5+5dYXhe9W1eAOE9HF4eZdrRd77uftOqlULPTCE/0KC
2mFtY8NqkyzMdp3Zfn0x+UgNjwQqNcEvppB6QA4QVDYwL/MQKav9cH0jPlD8r5MT0/QrX9rKZJTm
zD9RZyifaAOkXZvlDUoQKQrkhEZe7hr7UyuS32kXqIMY3XmxW44zILE+/JHWio2VzYlKWiFGslYX
TyafxEL+VmFebPxWuA12gfSX7T7thmnknoFeypdoNrHaaK2eBe9ivYkjHqzDiDMHpxmTRZ9hfuD8
BnDnkx3ruVHj7FQFb79JekKAhkFIxESeUKVqTs46icsOQVA4NiZ/UvVne2vcp+hN5osCL2WG0ulX
KxNlVU1uu8Z52/MZx4iZV+X2f2Spd2LB3iRn/KrMjAHtC1lMervWI8B2/gRNl7udUlhsvPKfvJJk
ip0u/mAeXGJU3dNSCcZoDVj0tbowVnhtBHE06FarOwxm/FDl4pSaY3zVzqC6HuUpnt8YwMjAO85Z
E70nHQCE/N1IuDze46QuD4R6DaJZEQzDOJ6BTWCVvgkxuJGgglwFBuQ3ZW3+E0udDS2HuzSqpvZH
xEFO2jV6GTRMjIgSfOikQGGiNmpCBDpcJx0QEL4jsrdvsadJ5IPzHqcV/C9yigJasS/qusIIWWyw
8Uy/kX7DaQimoe2U+62Bjn+ugA7N2iRXyuvmNbiqRv5UlUWZrARE1rsnCnH42A/encz7L9vZyG2r
m5D0J2MGajv+S+RUGWxbRyPkNHVAmkW5823oP1mZ2ZbzvoYCIMG7qmQBOY/4RgyFV9GFd4uiShgj
5cnGb3GLYujgdBJv2KFXp3dAg7iULuJbKZqwzZZEcD3sFBjqASHMkJWY6s1WEnTLH+Pv3/5GEnKk
SuZWp1otyP50nYwJFUrOmzSlgju9wPprcB/DkjqD5xUm6R4owtCK2huzRy8V8DGWhsLozDjgX9vM
jVKTvoai+My1o7fvArc93Px2iz047/+C90bozqYKREc+526h0UV3r9qMTlBSuJlSM6didneUxq4N
C45tGz2UUBXjozLFsgy45UGoT9/J4Cf2iDeBAQ6GMFXpTHPrQ7vsZb5IBMzQjoYPXS3F8PUrbjuA
gkL9ERu3lOpoFnV3izDupAqimQj/9B4kMufZ6IvjEckSzmwRz4yCXiWfjKJZ9hMRb8azm9rfI2bF
0RUAw9ZGrjT/8FZ2dkbDnrDIyZwEn5GvY7WeyISjW/gn0q+aTFsf4a/4LmyPFAlwNO8xMz9thJRS
nYmGRiXE0Yy0BP1qEplpV0mhRzqAilU5YVfTIdildYm1/Q6/6xmlHWVSC6fCxtB6s56Wl2NtCPiN
c4m3dAfu1agHZJiQuHpbrtq9YYYLg559cV59YhnIZ1f5ftodvegZBFzcCxY83JdI8CCE+Z55mtSe
8H4i6H0RUcbuwiUz3JOZtuTk6JajK5YPx1DrRkgQQYuoI6a1JeH2c5S/HIkbsMz2oI3vd8JCNGHI
l7sjZKcV9W7fLhL86QtbzOeVaCKFnL+o+c3LFJB/m+hEjCtdskBO2pIAz5Yl8pixHXTl4W9zeysl
jnhjSD1RC0qW8Djh7TQGT6KDr9dt+iMLF65vOdX/8drT0c/SpSN5PUB0ScGTnze5PE5FNEDMNGB+
xLZZYaQbztMy4TKl3w9q92CQGWkpIQP/SnDJ7Q87g3WI/fQUwEjZLauf8+xhU6WznrmYZEcz6Nt8
EtqdJP98GuKE0bwYlT0wxam3fkDjD3iyZmD+eNXPHRYJY50/jy4lBQ9ZdhqObObzgmISVw9orRz3
xeMCLgbj6BC8b3AFfz71F8cHvl3TXC1lKoxcM6/VYGfpnNjSDKGkfFIcom8jyUgiYzZmlVlEdE06
rKlTL+WXAd0mkH+85dSXwg6VcQoPf6rrEc7RLTw+hPw5Bq0clPKUBIFJ2ynehmu4QF5G4uzH8fqu
+025Uy60/Pe6KnNXKHRKoELSS7TROmTSYT+AgPU0+KDyg98twhSblChLFukrCOLzpmugS9JOo9Cg
A33jBDQiLnu3LvZL9ziPem5CmghZ7rbyGHA14WlBmemu75m8OkGXTQVehFj2o8Ee1a8fYJ5dXpGR
BjH+LP39m6tDGcymbthGsWEdLQgMt6fzo/7/RkhP19tXsWdChZGrNHTL4XycumLXKeRJS4TQuWzj
um5OKDqN5d2M3IlETQj3vJP1RZ0uymq8VNMdKQ/MQyTfKRvXk3L/7bE954Dr1pjqubG7R0Qz2Nif
J67qUnDgvRQV4z3c4TBSsMQpQU8BCUDWT722P1MPxDs/B3KbupMyykf/Zlwf55/IPk8OqoPUfA3S
1iBbYmE7ZR2VmOMK4u5QGO8AXLLiP+HzmTTCrJdEH5VSJTig6P5hGlM7WdG3J/IADQOsi2LYAmCq
cZrryQP2GtO3ZlQ5k2o3sNoY9a3WpachO3bikxDnstoAuMiDo2FcwQxI+oWP6MRtJgYMvNHXz3Xd
t+/60rZtFyRuSXpsuUjT8R2HtfOZOQ4RUmjpXTQQQIMowmcwbQhUZ36NySOsi49KzM8IegUHFzRh
3jYaEQZ/znrTlTNRYu44yR5y99pF0JK4Z8VD4qWKFO5mpNlSRMmrd1L5E/reOw8Ho9Y1NuRJwuxi
edewPIB+1L5DlX8lNTqO1wgdb2/EVveN7ruCAv8oaiJ7KLNuC2F2rn/WRRGM07J0Z8xLxzQ4t4Df
dhA0XSvj7UdTCAX1z3UKeCLSv0oujfjmfVxSkPSPCZBRo2Vf7uCdn52yHSzhw1C8KkUUFIOjkZFa
LJPmMXbyGbBowtS394dZifixW3bFbBq+EcZxalGZzZ2x4FpZt2cBIEmvX4c3iyMd4pBbpnPfKgAW
ROGv5dl4KTLr2G5QLW9Oay1eQaT0qSPiZZltEKOtqnGQsn3CUlp9VjzhiLzDEhYlJ+WKtx5DUlv+
IO7aWn4WW3bSibHmdEqR3xiRq48UmUV2uV1c8TTc32LTrZJqTuncCxMy7YAIGHSDM+IjHAC9vYDx
73fI7MUDxSma0yMVTtLI0beKYks8g5wvg1/KjV7ANWfrZfHaIFZUXHBy+tsXjiMtJU8VqT+jXmCq
26ieJ8KcE3LK9JZ93a+6BTpLukkGimVJ6nyhNO0ccY6SNcvenxukRSq2iKwggQEfiN0CrXCqSlWe
XGeo0QBhU3i/8b2YWYdbwJNaNVsqIabSoBYzqjseIlayDldfzBzySfd+TT0gAuD9eW4jbbnflSuP
ReZkANHRHlqX1tDCKt+3elBVfZQftCXUg4cw0ow23Us8fqnKXPDeOkSWGPSmKppnp22PKz4sCgb4
FxsDpW9dwNVkAxPhp8ugC/CIppM3N9Wxrf7u9GUBW/wI8I2pfl4KfXlQqvXMZVOTOW/GoO98nFlZ
JieHGp9osuiM4+rRFvI45b8NMmjqhdaJZTfI+IimLTv18hUdYZVLrCJGW9SbleXjPUBv2LpPJlVq
ZDoIZB8Uw2zdUgS4z1frL+Srbkd/SqD2tfb4UdnuJ/h+ORhG6yqI7T22g04WLBncVuH0RNXeSh6N
lA3bpe68Sw9oUDzWo2ShqMycuGuQ9ZnHNgQLUR/NCjJwGYdqpcGJU5kotkoagFQ3YXvnXi+Y/8/y
T9Vy9lYzv/ZOyUuKKqj3YIEnAY5HVO8wOcCm9VzSYphPnfDu2gGEI9N7F9jhnfbwhz7NY0txnIR8
uri3GCoE8JaQsFw9i4WZYI9sAFDZEazuRfSeTW1fBeOgOBISCvhstrMutTQp3aT9+KPl/dSKlYCZ
XW/0FzDQPm0bDgcKA2C6FFPFONkjK2lrx0aRdMpbU3vfjSIHATOcR3qXNV6+Y0l19R7jConaXNyx
4TWyA+4HsegLISrxjZq/Fzcofqr/420o1J0JO+6/ZueNg3AtzgzYXJO2bIvkmHqaRnMF4ZSiEP7z
RRv1iG8fyJfo6h3oBHDbUi8WPIQ2OrIxtrN8ivGf/nVtKgIwWBK/ukjuF1faOwZcpaOPQK6+YQ9/
4OuuDniMpV8FCB/xzLPHsaSNPu0NlqrrqOCMMBS+3SsreTuJWj/ddTAc4yb8vT9z5XhlQE9cF8Zj
ZCvQhSmZcy907t1/pI09/zbgCktHt0kMqpYS10b64kLnZByGLsgIkn6/3HuyZL+ytpPDKYErj6G5
WwUYgKQ6+mKnYUGqBkrcy2K+kQYgZg6WnaZ3neKSuAioS/UVi35GEX99IlqAbIGWCdNHgdi2wxE9
UGd+lvb4lr3ulOjEEJpZIQK9JSNJSicMnEkXtacgGMrnkC3qTGtjNNLLhEmHMbojikRmdvsZsEd2
8e9DyResxzcRhyaCTPRlEMG/ELKLEGOTSKNKqy4oCzC3IUem+lKwE97ZUG7Kta60uPQjI5uxx/Xq
FslEXNFcL1F+oSqtASgIqOZhBe1/TdX0NT4buczvofL0E7vgkGVB9nEjpw6UyFBNaads+iF0Lb0c
9KnWj0ffpq3pjnC0hxwtiB6RIsNZCrARWRdlrb2p/4W1KJ8Euqqm/4l1XnFumdlRLS4l7TxZj3sx
ChlAnnuYgPx7lnmg1W8Wm/WKGB2GlUZ1eq/fGC+eGnJ7qXgsGEdiUBORrpWETpE+GGKLFkALIfuN
EgBJs16q7lWxn8YZvNfufIyv/PkNaEj6wRvb/yiTBTJCVZJmedDareub1huUQ3GkHzGTbDygxpFT
/5WYATlSnh9KlIDt7i1dU7yUenWfEMGvDFcYC4JKrt72jbCibq63IJD3Py7cBDqARX9/TN2NfnIE
3UZrYNJUji9o+2LxP77XqjVOPDAkJTe59wC2tOslq1OtvW7NBOiEDAPYERXqrRxx8Lut6GhNhFYf
KR5mO3HJDVv2PNbRdV+YNYFRElvjzJRJ6rusamviMVXmsDfTK5jMpjY0/3ZK+IyGvfPO0S2j/gCk
iGIwhB0zVW9OURUnlbCNzzH+ZgaYvD6gxX1UlmfhG3c7tlxrczo2uKvtS9JhiVF5wB4NuTCMFLUb
B49jbFmGoPs3C9PGpGtJbnO4LiLoxQtwGoVucYrI9Qzq6thzyBEuJeOVfzKMxJIku0fwLj3LRjgB
Jt1Qej54xx74TMEZfO+4UocQ9ayqIy9pUShSJMxI7XIYXG/KVozKRopq47TxnfRaGJKIkIpGetFr
ZBFb6dF1eH3LD6Q8oQJVsCjrNJ4qPocyPcf7zqoIzCceJSWkF3RhIR51pJn9KBfYKkOgykxCP2OI
+1JxWXmlWJ0Q21TBHdvi6v6EBjeCOh8mRBPbtoUX5RyMC+7kEJb3xfiJ+rmqBq9l9E0PiDejWTmb
4MbCORFomyTSaAdRJUTMvXjOPl3yDVjgwBB1b78TSXlDUpFItOtZePw3KcVSDTMzqrCzkWqKRDyD
aMFUTgpCK7eL9yRHkyphtEs5EIOcbhp2ky+Hu0odTCGqVZLzPh3nfSQgyjk/IZNjzsimKsVYQRER
O8XvA89AvyT5DQfsHm+/0UrMhIN2tNiatDSYzyVctHL31gsGygxCJkvEQAp+Ra6048Nr7+9H4gJ1
5nNg0/8cKpeDLxI9wnaI9mKFBuz0pPJ/tAJX2sSzI53GK+GiGEQ+caMDTFjzKnlM1naW8OhWfHlk
swTkLJkkEndn4li1wgdPJmsVzIRSn6KR1Mp/F2H3/MsWrXQMFohDrd2Th7jheIw4gUq5aJNiXrTC
6wryrG0b/UOxq0ubUnBDp6pGt9tAHZ7FbWH1FUQZHFagAZ2Zt9YP62dxXKlHonFbO+L+qQoDhJXr
lzm6Cbz4YbqKmH0WGKKW3ZKdOGTg9KYzniXreBoiQrLIMOeU29n6q78Yu0qEJifLVe6r37+J+9eE
fNc8r0n+qk7DHA0FcDbz/l5ebXY5IQIRoy2G5kYYB4zyn7FIIGySxDJZk3fXbLajwG+dlqbE3qnZ
U4m1qjkBz+elCDWhSywt5vLk8DqVqbQH8KRJ5Vyj2V0ZH08ZWEaLu8LUP0sJxIoCpajkRPhFS9Qe
3sz6me/hEhIMm40eI6/K+2fSqpnL4jBX5pBAOiT7FRxnNoKeRRGsbnmVYDxEeoqBjHndIqaJCRsi
61QcF8j8giZJcHl3CUfnnjDExNX9dLa5lX8tTIv4amcRjcO0OiByS4YGxgWQQfnfyDb8Zz6RPw/y
ivv+LcgL0sIrw3HlwW9H1NjvPoI5qcjGA1vRoHpFTKywMgpWMPHDlQx2BXMG9DYevvcM5Af4dJC/
9U3fHNUMFZqy5afqBdLKm1xFZuCvuhhSu1xW3r2/pQ6X/ztEBc1WdW3CsCMKQvH9hmzr8Wpp/LRJ
WAVklBzsfcqJRzeSTRilz0iK3JfqFpu4JDFeAWaKEHN6SdkR1bqED5ueeDgyFLyz/A6M1jkkwfWC
PK6IoWViZL4L4PAQ+7EgK6NFXvcVxyxW0x8gk/P2rwmxS7bAlSVJdKRTu5E63XALgs2rQY+SsUB1
yleBblst8/ZFaIgvJVit/h1acJtHzm8WgOEZSxU56Zi6KjKGnI2PgxopWV/wJKVR6mlnUULLX2T8
X9uAb1VPmXr8M2znUdOKIXUCcb7QzoNIGAi1QHJJzE8afSQbAhIJtAFaCq7zUQEc1ncSXa8oAaYK
Jq+hHepQExD4tsxveBXqzbD6qRnHAuDd4udWI+SXj9jvqS3q1gBn9r+m+eJY33gZRkaqrjN4xGfK
7sIWTZR7jgs1OpUYfQwNpiJa1fMriK5XR2sDZ/pvHjW0QJibLwe00B7bceWpBJ5vT3L86oz75Fks
yf4YBfsnfRtuYcF27oUk/3Wksyssyv0PEOkF7g6gyc3n4QjyRg9pGxUg8GR1ez07RnhVrYUOO9Me
6zOOQ/seamzMPf4nH/NzulhCvsk+pEryXgPaLw5oG7ehbCIC13AKbBjYwCzwJ0noyODzqTpzb9e9
xQsGxMgIxlvIBb9dUKhw+dwrZOfMrSNEb8eYcQj+zKWAQyFtxAmb0ijA/O1g61wDxQUrzLbaUrIl
ZoYtOub9aLdJWlODU8+aURucrldPQbL4ba7ATEKLQl0KkKxb8CvpX0waPvdWPqV2kyiSHYe6p8zP
EjJJtKMxLOvQ00KYxtkuA/XnvX6ZqEEoMKvFFhTEaOILo/zkBJi7BB3gs9lnX1GtWhBL16UJoUYh
dFvoHzHzq5sUoob5cnxUFSdyLHpoBegIPKqs5Q4LhAuNv2xgFBfFsW6eAUqAw7oYd+N6JBdnKK27
2HPRdLRfz9rBGRqSY/qa8RzC/QOSw0BaAfZNGYq9pWKbdni6l/sbyHXYQ+TZdy5P3qsBV78f6ct2
+CGAwhAvTLUtM4wbRKWsjOcxeGCQgLPzznvJj5rVIgtlD4COUQ9JrzOr8L8zmXEhToYluQw8o3Rm
wUZy/SylMWlcT0jZBeSfZAAMbqqhWQdMyN+nFpS422AAv/bvliEYYJazp+xFJ4E4lKn95ftYpfEv
OihiYeGvPYXfOcbodAub1PP783qT55PMe2DV2sbGVJoKjucmiO1i5OgrSQKeYiCl2ITPD1evzdxo
yrCI4z+qQ4R4CZmvVbjozHBQurC6HVhgnQY+DU/rQVBGasQJ8F4RDEc7keq4u6WkUtKsUFQzlrLh
vhY0juBbFMvUzrFgt2rmPAESPD42sEaeo+zmlbeunt6uLbc6RoI48CrglAdQAqC5D24ALQ4rkU/H
NkrEilwwnrxQV5QNSK9DqDvG03a30bqTbHjznD3uQaTqXJyqwrvETrIkYoRdorwgINYMAD4kbury
+QpgiY4Q8dsLj2Qo0vtP2Hha8Hq0UUwcpZTQX5Gjo564g/TRwNvqqe0qvrkV5anvM7n+KefkeLoK
Wv2+FjmQ6M6yzauWvpNrjlHqjGbq3QB5mAi33tDX5SrbM0p0j+Nw6inkfqqhlP6RqpjaySsxRNVN
dj3a5kGldge2xthJlBIDFDNkMPAUDAQFqkTyDiboA39jlaNo136TNmhhyIWvICJsh9fdS58vLa2c
kdrQc26Ia4sn/OD04mGlrh6D8hAQQiCZbFup+e44x+PJQwXa2b6NXw646L2OOxWswFgJX+/VQdWz
v7sUM7r7M55bl09NQDopOYScbLijjP5VPhLEHTPrZujtj7UZJXVx/nLWegRqIetAJXiEsHvDRRzK
Mk84YYuF0bU+YDuW0h+D2jImcLeWeMeSeZVj2Ud51FMvvD1CpAV0lis7XQoaEtcxJss1PUzgMjtS
ifpEa/Jg/+rxgyxRmQgfFNSp6DJ9Q1kmTT0NaO49OBBrMUiaewQ5u/MZNpYuRoyaEJ/bbfoTpihJ
xkeHClIBj8CHil6uydQys8TrKdKKkVJNtUhBI93+vk3f3nogn/8QAFKxwgrrOMyQXDU2Ubmu8rm5
DJBROAVK2Ek+63xBeK5EQk6o1hxChmh0HYrmSftLyvQbZ5raSAY2BJnjH53UlRNHT8JHYai9QBDm
eBzpKq2LywZ+iRc2wbCA4oJovrLqdftgXrpole8SUxfDYHbCEmZnUFlbU7wCKN4zPpG/8/f+8aDV
KamLd+wNatyZphM+UqtRub0tNd4aFyg+ytjJHwZ0ytYTJjN8QdHRW2Apn4igtZIRtTpOggBlAcpJ
fEOhVOual+r3Si7iVDx9MAlFoMsZIP88lky7RCuD8Nr7QE2+UQLGZaUwrdOaKPQ3Npse6Lq6AQ0S
E87tsQRsOLSlAah2s+4H4U1qMHTyLpb3b0/UZwJXaVes03gvli55eocPGTZxpQKIiH3sjbM+SHi2
nU+ihc2IlUFUKY40oEmwEYcit0vn6fva9Spt/ZKcnx+NXUSiZ5uHLou+MTjHgCw5yY8WMBDeEGhE
MLCNZzGg87MGUer2MXRgvYV/owJrUoCX9EYLXlkm0PkWNpJLBvmkyG5N6bxq7ZE4JCsp+rLHjYdc
bxNAiwUf/xodZL8uLsM4FnKzchQq/MPhrbkPUSZH+Z0zqvR7+OdHJI3+IowHVjoY0eJMPATwaN/t
CcL3JpiguzKJNLeCfZQ6oeFuYPNEC73MdvcpHR4j7FbmNEKH9/iLSjT9JTpz3DQHZ0ZFVDAnuGvn
iGlmBK3I6rAtHwoywZsx5Q1zIoB2PlR7pZHPu0LvGxYBguDqcwxwOz8sZOYg4ZIpc3XLke6geyge
BSlofP43iqPIQ5xrgNset+Cw0nIrwK9lItFmdpAEofqbp8URLyAcPlx+fkbgoMKMWZapidf3DIXE
E+r/Fu6aJtihcz3GcjzvW2D9AgBMuqY2zEXGqSIGze+ISH80J6fOnONmInjcXORMRa768VWeQsb5
1sQYjXJOpEkm/+mqxvrqJO2Y9LBkJhEeIpyvFhuFGtfu/eCW7VNhYgO3FgVElEQlwgOzZtsaWcrD
nNdxInC4Hepz/wur1k8aXQJto7Ie/fz6Lg++fJE+Ns7823g2rIT/GkDr7jpLh5uFlKjCUsKFLUAe
fOCcy4AD/vLyD7u84nbUCsNTD+HdZ19aTtoonKTkRCaAYRSSdUtS3y8JS0QSBWaSmseVuMhWurg9
AdnZ408qkk35bxjWD/ZGNXz0RaZwr0krpmexQJYda13BSFy+CQXOGf1sJanuTxFA4GSLxxem1xSo
k1YegINFWBeQYcVoyXEc8l55Lr79EaVaFhAxnEWxRer7iKTmBAD3u1+SDKsqTMHImIAFAn3skdg+
elF/EIPHnlhNjsdIXvIxyx4LPxMXDNGYzE6GrbXQlWMes+OLBAi0Tts5S4XD5VMN2fCrRJQa0uA9
y7KK77M0AiSmFtihG10JI1zjexrMn0sVOfaBjvjj+D2FH34mbacnQ9dRyQBIqUWONXLRgQcfYvBK
KMgr2vDohtfUPrWY+eLyXrFvskrk+JXyasu86lY+IDniDWoHNGNiWPcAhgLSa/wxh/Idzg/hjCWw
TWIXcmJWFgzaCjduTXHKiXg7BNyNGmSVh+RV9csB2Np9nVoYqAC2e0Amn0ZD/JG/8hIXszOp+HBV
H5R9mH9JSoMNJz/TCz6SkHSMbtw/Ea7Q9BkB6Y4yToQwfupJTPNGGQ0pJ7LIbEybeyu6EQTNjimw
8v5ropBuheAiO18Yd2ikEOlLHg93IUZUREPY86U53bMYYYaIdIuRdUT69XDyVw3KnkoNNbuZvQK+
549ciDw9hdIojphjWjp+ACPFD1ilACUh3HbYJ4kKnsAMnyzomX2FoPbyCcN+Esc2pfFtWyXvOyhw
9Rvlz/HJMbxMITB3SeFXw5qWKxt/keLR1mmz+YhPkrYiCe16zIp++hNAZPMFUOS4Lzo+9RZ9Qs9x
465RyA0n5YZNJXlGmZDBX+o0o8KPQhMTZf6rUrOKD83sOw3PByS3VUs4Kf85muhBhTmUIK2Y9qhj
A4f/RirJDmIxO8LA5fLL8LJ5Eg2siP7MZ45o8DEOSFmPlOFZgUC+XC7YXuO/gEt9x1ketOs0QYES
Mnotx8RMv+FJgsWMsSv6Yo9US1mRIAHBrZWoFrr7hGRxK1kfuvqynHxUZ6XsMX1aQb3IeF/y+SIR
5VMYZ0WErcIzKdAhDnbasrixd1L/vKEaCJVhRN5JnAMFYeuSsAnwQ+SNPSAUSXdiF649nDeMKBnK
k+yfNpKlxwmdDubPtDvwQrGkhekSHNSG7DawqmEvjYHSJkfhFt1d/a24Q0BhfMSGNh6daQSniSRG
kbmlVI+lmZwb77ihOKWA7dKQl0e/jptOnS7IqUz5b7xqNL1FZLJ48mCqAi/0D47pD7C90+V7d2rn
7VpAa7JqLz1/oZhBvljIGPlIgWEM30hGC/tut3O3mQeCD5B/Z3mKOIvMQqaQDwQNDhq7Pb08GgFb
BkA+fHUosUtzSERK6JWUnVkf6ycp4StqMxbZHpWhyEBV4QLhPtb7RkRuo90YoXcZbHPj1qs1gmcY
Amb7OU8L7vxtpVhWXzQgHFxyW7EcEP0GVo5yyO7d2evj5ArG18EUXoHkHfGhbeRz9WpAov4j1FWH
BgnSBdZ8GHaPR7qXS8R7nGFWIBkkLe83mCH8Udg7a9T9/4eFPVBfMP98YZUY/BmlhXZSO0oQhFa+
De4+kBPDMMKBu/r8HhnfiLyzHAitxdTWu8ifxIdIUhHeg+eJ56XQFHbbHy1uQmGdClLsc0cotPi7
oIW4rfhinWzco7cPmKE90CEZ7VITJZoWOrMQIw8pjQo3Nb0EFCuFhCv9u+VOxwp61TkV60wEWQI9
I9TJEeRhstUDfE0x7EiPqmC5dCLqdtKYjHi+VRysczCdEYLhyVgoUg0az0W66TmnZjR5xp+kSjXw
AlC6HqMtHGbOSJ+oaD6A4SX3NiPjGaMR3dyplZUZGVES5c1ryd1SfBMtCm/VKfVhSfQ6K8Majv4X
tPdjpYn0MEzUBs1Sb7JyyDlXyb0fSX5bhoyeDqEINXxBWpfjhV83Gl1H0OMHGYiWaYVjyU8dF8o5
QPdbPdUcsriYQMCDLhlFb9xBZb6zyrafCkklfooBi57cP3NuBk0dmFBS27fuufwhwTHJrSkp+dmE
5wBsfkjhH8wNsY2DWI8cxhVjc2UEvIrHc0IrBh0nCHAWziCPhc1jIPLAcOGTqb+rIkKsdqXpWBmQ
mLbO+6ou4Mfh8u/lyyWVwxm+HLtvJCP3Gsbw9hbE0sRhgmSKW4x7N4bteEhGx04rM9bTUumnyfcK
VeZIYXcD+xX0WgytoKDY0hyLwYvKgWu2JUCywWmYpQCF3CtmNw4DMddXA41lJeW5r0pq966O/90A
vSidnTdPTTBWLRukVc/7XCA/a3n7gKBSicJsOUfeqdCZo5nH9YkjCvqyPknOll/xvLGvmBRfsd06
L+ZZ3o9l3HttLMlm+/h2SOr3xZ5OE16xoV23zdewO8UvTHePGRpfBTZX7Sw3tKN9mVOJIeqKbz01
oV70eiqAv5U4l3CLfVpOBlJc+KuDg5/DBd++spnamcbWm2+aXTKODuPJgntbn2Ro2qn3r66kZEhk
Vf1Xf7hC0KYfMsU4PG6UBT+/Xpllh+i6OU/oaGwse+ElRgcOP4R3CirnGIqiGK/CdKc7NZWHyoR/
POimrjhx2cDDPRmZeWA7+exvbW3I2qL5qSql4ZM2GLd38zh67MS1G5S8vk5IHnyqkc/gPDz8wZGU
nS+bQINqWrKGUbCXK47I2f7RbDsfmfOxpGlbCzT2NIV2yra2WEv+ZhxqCdUInZHNvYv3gzZVOPXo
OOUaTjsaCzZLuWvTQwtyKazBLYv4uGxbuVJKgRRa2k5ut1iNtfFDtZP/k2oYf8/EEP30zURq5Uus
c0bV9JUx10yapwD9fmn18Vv1lEyOns65f2Bd9oL+XEao6OUlesljwTFK2WytqTZUrvQgsM7epJPR
rYRzPqCdkEF2dl+UKc3kHkgCfhrllqSxXslsGyrfxssEGxuvDz0vybbR5FALlrLLQD8di5+PPlMO
dxYcrviYG4pwKg4v/z2pQ/3kbo19Q9fp6dM+dSZR1jbKXL+M3frDa8mtY/k0TcCEjPDHlGNQ8gzv
kD9baj4tTmZsVyQ1bHqC1rq6dRa/NgL5VVdzLaDW6cnnUuykUd9mlWzhcASMGabf1lFq1qntx2ld
G/qO1trsIXVth/AiVJJHtz3pYAiaNpJzf18J2DUc5u+J3Z/pEN/r0aKW7uCvKaa0Vzsx/TZke14H
U7RJZYu8lqyJ50M8icVjWpJDdVBnX976YkopTNQiNiqmqwzHepI+OVvKvo1LCI5xgtfLVhQ6LxyW
dKLYaUtfMIrDv2onFgGYPCZiIiAdtPi+5RKZmuPNmbIJUZiz5O/jdLbzHePeb71n1TSUFre+xYSc
0fW//j/jlNxwRmv2Zk/S3MahKGRR7uRLKlYaroozLMLY9IVnSyl0zQEJhGb9BAFGXNZgEpEVEpfz
EW56Bf3i8xQeJsXaWTVROBH7Xg6PYTIUXMiJXSs+D5XAWWqd9btLnWp0yw0Wc/+PXlY8mm7lI312
U4Y7u8OdnBlJ9EsvAzb5ERicu5p45b7jxVnpgoTYvpzY+IXoOoQqRXGwjwbx8vKBPkqrmJ9mvnkN
zH485YmiDDvoX458JbFDTX/71I+86CPSeN5MfwgleS8lvQVY6EHJJm3IpsVCkMN9ZBPPZk+D56HT
69NMVBupSKPWJVkqoyVHuufOgXJw8/wRrXxBv949AnheotmWsqD23dwdB6mcJNq4mSRYq7oxCj05
ZZncGkh6LOfIeWguJMKOVXajUd6E3wCJvBXWDraAyIKp9sIUcnwW/ebyU5OPrrAbd2/Yeq1rxnNB
2R3vjY3QJcu4fd49cFBMrpmXwXgo0ERUu0V7KAjcTdzi1zoGwli6RlseOQyeBB/xBlP6ZSO3fczR
KuSybOLqiOX95x1SwzCGcpTIJPJ8N9I0PFe8l7O+36rwKQs21cpKta5RqdSOsVb8FTGiVVrlxrVq
gDlUBLPq824JZCs6xsS6VPlFOUWJ+nQYW1Yh6wlhlv9exqtWyZM8SCTZAggJnXzwZEk4KHBdXBXe
mT4qdCzkytUVtxze0en8yEasdMySuc8YnUPwQmBU5uHsC5IHKtUENh0/hAA4EjLSAS1UbzpvEprf
did1d9HldVljk1y6ubRnz1s4LlueN2BjiIWYEGZF54yr7jOMEd3XcoQkmhuA4LWvHwYNkq+RNYWu
eyya11Jp8QARo2F/cwEF/MvQw3hjLDrdQyvELLUer1siVRlHGyuKT+8hJ88rPJYNqiWXZ3FseJHW
XM4+il5OdSkBsFQt9zthHec5sNtE9+gXM/HHL4TuuBRpJlWGctdWIhPc66G//iP7krgKoweussMo
uUXJQhuHI58OW9HCvsYKTkQJWf1YP/s++7QCbTv/rXM4QCLNcUWVYHJ+XUouo0/I98aLRVfTJ7I0
avKeyYL2IhNRJ3Hjh8SEe4HlVKUjEYIXlOLgYIvQnvVDCFfxOw8pfeoYWWcoSUwkRZxtJ9+qfVXc
XCukeB90WM+lhzghSrHfx95ppSFzs4bFuXiieej1Y2SChjXZOqx2oZAUy0bvr+UbjWomM95aE0Dy
g79AFfq0DfLxsZ+kMDvA9GQDo3H0+uYjdYo/o5zRZGar7dNF2j1SdtWwgZRRZjR7MoIpShKf7DIV
tj+O8fOECbe+f97oUBw2vuYOTPV9CYocx1UP6lLMl8r+EgL30EQyQIkJNbvs7vUylsVcvmnC+izZ
qXyId+UurSzzH09NGN8CSj92rDFrcVN0G4rZJKgnMvIK75ZmhlOkKc71ePdIjTr/WrBMB7rtn5ZT
RTISpS6PS+Rb7/nfit6cR7i28EHMMn9RmC3JBd20QUlsd7i4Mdwn9ZNP8AlegqAqUB8a2Xri6rBM
Ao6u0qaLiJbwkS7MJOpiSzdGDqjYKU25OvyCgDV/nFVk0sst8dvMRkSiySKb6i3VVCnYqRooO/wD
rk4aMBJzLIxc1TQicPsjEBTyfiLI7/+d5H8vsngCxF5thZYyMP8jTrX9/4YlUHp30eJW0RJjEyAg
IxhsprYA1Wqr0nfX2QKz9wOhb0Q/LUs1H+IfOatkzJGWuXbYg6B5AE+qMelsGgYIe0KD8DeYcsaN
bvxqieDTKaMxEIY0v+p6+aQkXcq88fpUhkRWIFYdiAw3zKJj/5I829j12j2gVi/dgDEqIMGuterT
UbD9gCoKi31ELl7O0GNCqnlEuSeH37K1MGqYMRce7WRCr0buRM4qSQs54EfoefTvFGcRJtPA6ptN
fLTRAioCHLyjctTUR4f3uRWtFfIebHuLdwIM31GEl97huDV3KIvPHgPjFlWey+CFNQhswszm6Vsd
Iprxh+EtuJSDFwlFnD2bI1g0ChVKR/5yI0CcERMP8xuGZv0yO234xRy/TqZKAAsXgV6ci3GNiKRH
OsZk826s2fqi/eQhs2QQlcBqZMz7Yr1MML0I73F6W0xhrIOePSfASNJ0uK9eyrz6w+iTLmP5WU9Z
YjG7uJdTTEUguj7kDxtpWLMyyECedRCORBWLjVdo6tFvTlnmS6OTBRFna8+mzJTAQuznCtom5kXN
jQ13mh3AeQpCuAP3lvWRTsfxIxM0/o6SlGb4SV58ydiExwc8+pvfduHkEXYKTaTV9YhdJHM5yTX8
Tk1BTgBGuEVu9NUrCiGNYM4y23RFhlTUrS0skO2dKiD4Z+BKxX5IkNmEs/8kU4IrJBvsR8yzQwFT
Xb2F4lmY+XElTsg/2zDWVQjPaOqWDKdxwkXIMyC46o9Rmo/F3JCBVhtD69BcujoJuYUe1c9+7Qqb
gZeiopqkOSJ617ONwu8tuaz43zktg9HGUzNXPQvILGTYfKT6r13qpEkyuJoEU4dAjRTVDJicKt/5
4aflxjxKNIgBy9qv9vgo//cC70dMf1KVkjzk9H2w906XxD3wp2zYvFNb+HmTaWdgXCmmWPjDGHKC
8nY0in7Sx2ThnOdrUPimrGvLrLaomYznOSBbqaDbPTFyhovJRxEgiL9WdUB9UE7S2+wUk68Slb2C
Dtr7i53R5KB300uj2tgD+A95BZ65qw/zkQz58S8UjKgOKijafOIN6dGtL/AqN32EE3eXx+jomA51
zrxGxu9okKvt/QAgOaqGtwMD197lsoydEzJeOUs1UbfdT9khPTWiwiJdvQs46/K6v0cFEtVqKMIL
cT+B6bGc3BVWGqArNs8GLJDQ0QYDkLQKjxG21QAHnTcBwVazoJmK90dr1cVGbx9H4y17jnEn8IPj
T32gimCj8PZ6MbUP/OrsWzscavcOXXjThwBed19J7yZMNjjZ+zVPuQmaIZLgDpvlomgrOpqbrcja
QWljnKZ2A/VOx0JbC1XK+Q9uFPwv5ydRoA1H478hlCLpiCdSIm72gm+jUWfK/T7IIu9Bzxs630Gk
W2cisvuLCvyjPh5+U1Ofhpvnz0gHDRWnV/O6n1Oa2+x2Dr6Tj6o3EH7/B7pcREqlsIjHgLUM0z2w
SsPCpqV21imyy00UvDojyV4RsGfKP8NKfY5lN+/bYYw7kXUNkOxhH4Vw75sB/dwSpTaz4mXcYAK1
+7+BYzZ9Nd6J7SXKOQBrs8ARfMLdEjvQepNP1dy5IfUQaPTB430X5Yns9xMUKMINcbNfd1bRmcE1
OzLbIkaK5dQ631LPhvB11NWRuEFxuMbMJz7fSyD7c/SdpjBKGzjbsL1hhSlUiPnng0vkS3TLvggA
SfRX5xxwxFR1/H6olsyVRAvaxKOwrjhZypkNTS1Y8TumrRG+wZle1I1qqfOML6dcT378m1+wsP2L
Lx6xL/2F/0BBtOcfXrA6Q6VH3HxzBrP0cqXUrdeFiHpsNpHzNzy55l8nb1GbhSQKDEomBXZ0h+WJ
bA9skKS3Ubrijj7HQYJjhG9IwJXYMFwD382w0ERfMyfWa8gCHxt9SqREaxFJRDt/K/t7CoEmimoS
eY4qfUNcgOYN68GV6WeRiOz5YERxAW2vpTyeJcYMvUvx23xH4O1IjZ+imQVC8Cx4voNoR04tHfpg
zX+k7ny5DRsSI+7nShYip3vuPFn/jYyU+6ABW+pCp+X2a8PpuEIrMdWJHSEDYvhB0jm0D25rq942
7CeACvB7HytmKXoTzjRyN6rrCT7dabO1DNWereH7kJ75CTeQA5T6I4M+eJXN5qaVdtd542y38N1R
qNMAep5Cibi5L9MBb14CDjXOU83YbUAsMdu1CLHa6/HsxWDzQ26HqdZ7e2bkzHuV/Q7iLyM91uvg
n5wHxqFAirscIuvwALqH5+7U6WzBpOCBYjX22N//ULlXrloEqxvQwUDL2GAZ27gMLUAkupns+ti0
yn5BkfJ/V9IGCEfCy3MKx2q+OdF2JMlHt79Q5ThvncsHDUPyN8HLiEthjrc6CFjTyHutTISz1u19
226vXaalAHtb7kMjed/rHJRys5apJmK56OrRfA1/QhkOTnN7HosUUPECbs9OjLlyhGx1uCQW7/d7
VgoYEfwUQQvxxoA7/sREBmJb3FrPNXY5Zf99mPHHXYpaYvpDiFnujCyUgFFAAtv3juAfHeigkdAT
kCu8L2kglwtpYDBHO9lVStqT+xSdfkoClvWU5dsWUUmnpsrjJA1S4A+NhmBg2GD/EI1L8rfqzYYz
qtreB5gqX9DMyB6ODA3N4xTe5aYIx9j5rwPAI3Xh118PDOIEDJ6e1UUwuvhNeTnuYo3WixOajlxM
Y1RvSY9Mn+TEzedVaZegO+YbHqV8qS49GTXkJEmKEs3HgwOaI0lHjSXqBbRFeV0HJGYZ2OITcY2n
AevzKQyKPSnct4DF0bbBc0s1hQxlXExqBqkH22dxNei9uIEgpIuviRAEnOFmySPVp7YX2czHGPYW
pqqgrx2EfbuKjTMQBS3trC0TKWjmjWkMorJ6WuTYJYbK+nu3lU+XGQnIF//C+TYn6HlrLbtyrR+G
vt2T6X2WHw8aF8/w3ssoAPP+6cdV9CGL9uRPa79oD09KLFaBgbiUaE6lR0CB2CBR+cBtgY2iSrmr
xbmmqlUZi1p43ghMmR9Ev2FpunkjBMC58hwNJdbml7kPf600A4GDVGcsn07Ua5miZkOMlqiEWgXT
55FoWHAiYIGDzH6uQRTAAG+DO63eWymfWpeK5tSpjmX/VZ7jCqkzHpnmDnymTgaObphCQZZCh0rj
BRFpFFlQ9Mk06y0DK/tSM86bEQp0oDN0BJxgWtD8a3d/K28hdnsHukjbe4IlCFiL4xJ4PztU7iMY
n693gCZ6kqiyjaUlUhFHoOHylUiFrYC7r43N4gsc7df9dCZ57dD3jiJ7EKH8gZyqpZ1WxLDa/ffy
OCHrr+3/Zxtd2R3hbbJ2bgXsUkfZIsngo/Yf16XxErLcijdB3ghOdN4yRwzEsOhos2ft68jiNpIm
DhOyil5qnDTovkwNWBEdvLLciY0DY3rTFqX1akQWpH/TbMwTISer+90qEBngvyCXmtBZrrWsyjf7
aTN3FSaGG2G7nEts5XhzBsa90lfB1GT1nGhwKJ5ZZkHTjt9gVIzzhvhL/cVRbaAEWSQAfDMKqFMk
DyPY6OvxNDdkhCsm8MnyIoNQEZdSM1nvE4tgAksm4K6JTZ5Zbq2dsNxKs7bTjzqz3OymjW0urztv
zcuSDx+aKOT2pTPk7l1niv/n6YCHR87IvaT1Lmc3T3kA0p8Ypa5IgzDyUezVq6RJxAIeOR4wFkyd
xX1Otc+wTCHNxjOyJV2PMeZtKTrV1fuwzuYJyB3K4NVcskDRDzoKT/EMEvF7tY0zbQKDmcyQVlcG
mXWi9CSrZsR73UwxpznZsEsL+O6MepEZNXAMJJj+zuY1lAbWrLOPRlcROR93SC7y/JRAv8U/u+Bk
3cNMT9WLiOfg2nv/CZBveu1qWj0r8OQSQZsABRj9jUeYcjJfhpDiMAxilaleqx9cYps04Daw3ySU
ijy0ZU/7frQATnwlFIvVANqQwl5jtPi/UokopqpxCMC6xiMss4/7OtFfozyZ6lRi4GLZFRmisXxJ
MFJ3mu7ZNMBvBJTf320nhIjauYDtiZBqC2kzWHSVlfcbcmleXHLDVNUrHMJUDj39Q7zT+iA2WmY6
Eato5NacAxh++4VmMqDp2ayp0AO0mMtwrZRzWk5F95tAC5VQCudVXP5GIMVQDY76CDDYyxMHmHji
mSkUZgrkh1ktImKdz4aMbqN2yhGbLNDpvlsLktD8bBum95xxdkaW7HqBswxoJQxOT9YHJkSgWkD/
ccmNwx+NAkcut0KvahUjv0bI57xoZqP/jxSi1eZyYUIVXwaq9AKD8fqjIO1ap4LZBHdbXMkl6IXC
tH/+sf1hnGf+MIG2GslGvrKIK3EqwBWkCiLUTppMSOFDQn2f05GyikZxEQywNJIGF7P5gwdmnEgC
/5jcmBETrVfxL9GOjk3xU2UrSBNymbbZRbn+0eneK/gCzYIPG+p/9cqlduTJwrrzUGrCEFeGIQ8f
ndXq+3TT36ihM2nJX1xduQXDeZogSKG/LenKamGMNUYs653lMxo3I/OWJsFxgj4s5T5KU3EJ7o3+
mcD80yneOUPSirMEk1SOnDSaT1uxVGZl4XJM9AtIgDA7fZNyUaOmukAnPMtzvoFkvLsjgiV4uYYf
nzFTUwAX1p7Yzhu63kANowQ1+lRRLZ+YflHd1u+x3h2BHQRkrs7crxxHe6h/1K8gSgxYC41gNjvK
L+xfMExdt3FMJxd20KBIv+d31ULYGspU/qEYH+ijQY+hNGEtw+jhpmM/98ceUtb9uNT8f+iCI0KD
/tFoFAhyGNzEMTXmCWA9PGJNX+KAognsC6XIJjVfvnY3r4vL4jCjMRNd+/50iyYSyYa4Cb/vElUG
jyE5iEoH0p2p2j1WLutH87Aa61/tYDBMv7UQdLX1ZwGboN9Vqp6o3Ihpto1u4U8lEMTsZwoido6p
gTLpqKArpTPVtiK6MAct2y9WQLGwwaMLfGYCdX5u9mJzhIstPz9MdzBHWM+l+JMt4mtftE5r3xjN
QW2s0vhhsS5BuM/GszetUcTNLW0x+yz17re+K6fkvqbOUHFL5xCmG58VqG18369VdvfKQTRxju01
QXQ7RvTqBbY3j/Hi3Vzs5dtazHlL2GoXR6w9O+88jAT4ZOzsUKceppZr8F7U8Vq1RNPIh8iFwZd9
CtdR7AUmvgGdOw6+TUPCnvnJKlOlA7qEQhzHmf+0O9KjS2PHqaVKinVzPc3rxet35VIWW0po0MS3
P9Lpqssu6f6X562GybFUACqDT6fBy/FH8RbcNR97/X290Vj2uppP3B8clEsiWd9kD7/3bCRdXfn1
KBDX3VUeYU8e92eEBh9iCsyN3axrf3SGTylg+SEFKzI+0bB6sZkU+6PfcLMHa2gPbOJsyPv2kX+N
551pPXdOHHoHWIlZ2fcf8ALZUTj3xHyD5A+vV8DjKlEXDkC7Ybd3URiFNc61rBob9ZlaLsF9cpjR
YuQqgNGmAgsichjD3h44duwN+UQj4TkID1sxiCUy6cU8FjbgRWEWNp5BnLD8CWifJAppm7gyM/oW
kNO4BQzeGolgmNfnprdrylAtRGKl5qDaM5iFzyOfXSveuUyZwC5resLnep28rTTBZRci+QkA+PzZ
WZG3c5J3SVCEBKztXxEOZIQoCf7WDDCeA5pxeb3/Ef1nmCNNxgMUN10LsRkGTLMUPN/pvIjTO2mS
HjvFFoR+HfzI/emev3JT/HzXika/EtsWax75Q7mheZFTmH2mW2m43gN9D/rLuDC23uitn9CUKvYA
bK09eSGggRg9xwvIAXi3D2dSBfptKdv51yT15V6/0e+dSluP9FVo07L8QOjkddLEWcsXEx/RWs7r
3mv89WOJ9qqms7PlBA0VViFL16iSnliGTKe6shLe8Ipa6YVhtnOnIdmWhPOehy2xT6n1Wjyt0xFs
xzTrjaUVFbuqTDjYR8NLidb5mg/lxUip8lZZ1H1NUshZMAKk83cELxoYbFCT5xDdyI03P+6odvvO
N+1Tl2JL6dVhEl8BmFgJSlCTOI0LioPBawIA2n5Rqr3hRslmCd4hSlD4A5Vj2L9r+nJ64D4SDYv5
8b7WMUx1X4Au/1IPn5f7xXQBn7Tyck1TYhDEyQHCz3MIMxwfTEu1elIDB2el1iyFEGgysxbmfJb0
7J2GCKZIIChEJRu3/WK8S+xMuO+kwmGC/Tn+LMkB3EY2nz7ICHT65unpIgL7E1CAfAoghopuGTX6
s3QiwDW15ZHA9UpgYaipnamrKQUPShFPP1BHiWUkGgHJu1D1FbJ8rZZLNQbA4qjgIwxc24xwNv8r
h8H5itGGzNhifBVpRwCeCnZYstktQBunP9o/jJ+/KLMUB68Hqe5HJ5RvDURfq3F04ioHSF+xYiSa
4+VZRAbjwKnetuareDHYVql1JoISMm3AizE6dJJuvyeBSEm5yaiTO3+qsZVxvRb0uqxy1If3D/Jd
meDs9g9ogtB2ZFDHwSRUb7rzqoju0jO6ed77T1XH0pjoGrkp+Vw5nLEOrPjX9xXa1VGaU68O1GlH
5gcX8mXXFMPTEiZRpFzJs2MyqGu+m7jc2t/M9xMy7hF4rAXa7VxVDH18+aKU37OY9k+nvRKUyA5a
rLNrKmlB5+EL7/A+hjADIkRg+OD0ICeUc+SgrdS7XvAucwGormJf4oHN2c+a0kljfV/+Jn8hiPir
UfUux9J1Pdw3ylU94sgtFAV1TcUUGV2vRZhgi6qW5aacg92xkxDAdz3iJyuiOjcJVu4fvdz5cwBz
rDaAbc6oa1wno2JervohW1t/LfzmzvQRevD/cwIDddpcHRNfT3Uz1iq96RjtID4b/pF9F/zQmwYR
q59Oh+7+WTMK/jxaE1djXB9fGXc6NsxbkeluM6Ec5r1hs0I3ZRbdwjxuX8EcBgnDwHeiSGmuh/42
52mcTDSkN8OxQx6JlbTuo4VmM/uKTCoAVJVgiEuS6xlUmPWKbYF2kgqIAG3ON/epyAoNQYvsnxMK
+pRLkPIgDfNV4mM7v4xkpxahP9yDa3zNy6joUliC1wOw7n/nR51Xq3er0Zcg8TP4hSQioxCusnUs
z1SK/c+yzAnuu2+n0RHrhpgxl5/4DDZltK44+f74AqyWTRVaXDadueOGiaaokUWidvR/108AXNlk
ifOThyeYrfBKQi3rECfZd4J3bwC6jEJxZwhnH3XIA5zFqny7UhBn/jF4n32GOM9O2HATE7Le0iKY
sLqQLXT7iYpXztWwas68k62+EggEG7rJfKrSagDj4HmokipCyiU6gPh9Meu15SJvI7YYfHCRJr+a
HdB5ylUgKj5NvFv6nPWFMwobWt0hO6+M6/olVOtJkQjgkToyqoBTIlVNbWyksJOi5P/X55BoG8Vx
pUqXcLMGALKUaQC3dFUK7HSWHTO8nm1ckAlwmcjgvbHkxUdIk2XgITUOUX3UO+5JQJRyaHqP9YIx
P/PiO/Xf28qutkJ1wwl9jddUcT4+GegwqTx/waBkN+o0I+g8ECZ2/wB2KW2RPGonwL+2j9EOk3ez
FmDLtaA5LKpF1a4nYTqhEsn+n41gEnKx0NNlgRi/TPbF3IZ5kjuQ+v3tWljPH3o62gVvu1CpJ7CI
GOmCKH0uxGyzr/auyoCeuKadtltQO8fJnoBS7WvNw2DL4LBE7puvI2rnQV8fPmTSZOZq/LwFaCNu
1R2OEWxOZLz014m9VTYpDv6bIZtjCs+1QZIWjvvtJ32bzUYYSblQUXJyNHJQref/1m83ekd5yMfH
Ga00nNI8r3m6Iyn43zCZS94kEFYClhBMj409SPZoZJYIGrFFPNVmFMDCfeMwu4FSNhqQs6nWMh2J
zk+fzhFieX+NXhAjnHnaMF/toUVxOa0mOhZ7vP3XJfjyQduCkSmUPOqrOVouhocEtkIQEIoak9fR
UZsOMGwovs0edRF9opIYmzaEm+DjP5hzFlIOg2rTE41k4Jhsobhb81Xb7x1S2Pfv5jNmAB3NgEer
Edi/dX2dQO4ApaCUpRN/t+mTOejcZvQZ1rJ9Bs57ggIqBXX8NjwwgKAnVaDJiPiBL/oNZ+B53oBM
GRodunQbWhSip9qO6aFYkXGCg5k6f992kAv3ud5m3lrgZ92lpqnfBfLBwdMJVaKVRXAPhB2lcAma
MR4kh3dNnOHO3VLBKDt32gSokQUA9t92pnTFudEmCuTzLvfmyRLb3ODnLUa4A0Osr7oiYCwUnhZu
ohIOI/Dm31ZShY+EgVllH6Gp1/WAf5ZS8UQuzFFkagox3+m46uYY2vY0XD9sdNqxU3F8sRcQmVZX
nloE4susNCgYnbL3SczcRDxBuzT7jKUQYBfXg60JFH223ACZ61e4Dqho4XQCBnz4cc5kH9kOpOlz
JiPuuoBt8ETpIoTJSXvI8yPvohzk+F/+hVqSuhqsHCbNEyj9d8lT3uOMPHyC+TboPBl3z6eanQ3l
nrPN5sOaiplxFkrsubecjbgK1rx9FiFxyM3E5QOGU7TQKdWhTiZz1IRO/BErCs48EJrHpCDRBQxk
QWBPALBMJNGa3mDw02GvdVA6IfgJPN1sP2w80gv/T3SgvNNwApB2nK4CgCt+qqM3HuKwPDRJPcZR
NboqWrVsQ/xzZFZhw7cjaJQa6evdUf6H7wUMctLQsgNUc40JVZdPslOchbaygUh9K/aP1stx7st6
NgPyZBrF3qm4JzJ4VUuWEixywDdvkZ1w9wT6gmpb8YsdAN8Vm39nBsVDXLDbwnQrJKaQQlau/ZWy
l1KOPn/rI/E2LQpBVaLStoS6D4nmeNLQxNhFYnS4tZLCgiR+Ch+WVWmTddVO3mIBB+3YYfocSXZm
NeQLJVsj83pdIta+bZovNF6VIcjnfo/bEU7feayNt8BssufMHjzWHgGNE1gI8j2ah4j2YhaDFpaa
7mHcDUuoGY6278LICrc8V49ksnEUFtIL8uUEgkpQaSsJDBqqoBV9OojbV28YSXbR7anl5FOGT3K+
MKPF4kjV9SvkKuyj5U8q14zUbpb6gsD8vWk2jX+pA6R7sr/q7DwR+LLP673/ZtvE8OtcIVr+nAXc
alDYrVtv5sZozCLFMIYihMA6c1jt5zqP9cBcAvJWqMV0oMh7m7ATstDDakWjZ0I0FbFpxjFdMvOB
eH0U+viRkfg124Wm7zhoCdAuXe7hQi/z1Z/YaMDzo/+n1VPD+/EKHBenawIRCA6jJXmqf+LpkZAW
GNNojZEOoFQEOz4iN5Nj8zjaqsCugHVVD8IpcdmJEjHo7+OrwRyF3xzvRf33neH3oM3ludg/huSt
U/d1Vx2f55ijEi+0fKBZcU3l0MliU7Z5yd1FE0YNMIaHqDuvlOXEcCO/7ZiiqgsshLVlsA51dfeg
LcBalMY64Gqo9RnQIJ0o5PPDO5TkDG73lU0dwYo0hHpUofyLy9aminIrOQRdBBIE7/p2xrtRANyX
AhUtVXbMpfOjlj1zGssRm6DDTS5aZ5IrRXAuysNrughom4RWZH0nImeVAZuqpBRBB5WDAAZTfDZH
yZWzfGi+kvmnKWQxHXdNkB+M5VXGnK20ykmM4k4iElzv6OIZeRB4qxF241IpQgmflniVW6L6NSC6
pSUXyGgnadiS9GI4algGITKp0bx7BV02W1qZkGAJCnT7gpX3lpfdpP7QW8ENALzIsI0bue0DTITF
Q96PgXXsNe/lO12XPHHKxEElgyGQnkBo2i018av+oBKmeVW7deVYAOKsJlYBrYfkmM5FO0Bwp0RV
cSaZcmuW7RUAur1/ipnX7LxIiElCXPS5FytDrrzEbsFr6mksx0bDntHo3cUKlkWhAhJEUlbQ/aj7
ca03hCllDsDzasQthFvCpJBHVjcK3kXZRvnHNCi4YmlpAy3ZgMbpwKO6LMPf/EpXKFwYc9weK+wm
IHT7FgzXSiT8UKWf1fsbaqBiz/eyaq6KOVBIm72hs+UNu0Z10+DNEqMSedH+gnEhQ+WlEWifCX6j
5Qq5v/QGTnwrZ6RsH0MNFS++tiuY4FqDrSezgWLgACqZiex+l6/KMCzcSVT5/6G+l9taInzaw0S+
K/VBtVf8Q9ArXeMMQun3K23nzXN9N5p4XY5TD8k1Fui1PI9J0Uxt5pgXHJITV0P6za/Lt5Oc3m2S
2nB/e4jj+GlL9kCPPOUxeYRAIAwAjkMsUYgufDUkIB4I7/BnxnN9Fn8QATxCUuxlaSqUFm9mmYrQ
RQJByicQIpyTB6/ixZ2Wyy1YlhFmekMQ1wFjW2Shu26oB5fp0KVG3c/Eks7Sjv7kFa6zfL7GYGZK
rxhpxl8Wg1QQPjhKCUWCCk4DXInq8jfmlbQ52qpaa2QSvhDJI3l9G1sczXC33cHPR8vBzSEYklVD
GAa2A/9D9wrszWbMVTE+NZio1pe9JpWEjFjezMsvhdxCiIe8OLegWJQIIpR8i79ehyxC4N36jVa/
XXit9QHPF3O6dNzrZu9G+VvT5ROLRwpP7mm02/99jdDrAQ5OP6muE7q3Q8uYQMMQfBO1PtiZ6mTe
hNMH9xqqxP45Ax0tZkVPlWHnqUJ+R2X9TduYzMAOvbmaZEBhAttYOESjcXuAg8iLNvXHN/yKYUrX
Jmbpo02F7MvJe6PPT+m0zGK48a9rSVb071Z4omU/hOmfagWYqU3LYrhQnHg1vKFnHE5aHYmo/z3h
Zx7HtCIj8eEg4DsFpzrSH5XKcfMFP2ik7FdJQlNwkn6i8LdibPMn2YbYdLWsD04hbslSEokvZAYW
XQWHBIVH8EaYrIpHCnRnRAmDPYiysEAgDvqtu1wdJ8RA816MGAiGfc5u01GTwejYRbgYkqNHRkNP
RSp80a7j11mNrKYOD0j2dg1w8mV2VRQCEMk6HQri6gIJTCaLNvcPYpOHR0/a7H9ADYn2UnQdvOUu
hzdAQ8uLgE22JCXNPR0pEySgW83gW0IBrdD4K/F1DCbaV/Sk2p62T4276NXAx1xlU7evtjYRrgXE
WuRuu9FwjJi2g7m+7WTpCFnm3HlE3H1pV4c3SfUw0i+T404JlJ28gF/Edq+l3nRqaQSl96LHO2Da
fEGO31qL5YOMdd8A9NHHXqQwtAvrb44eVqIdjTK0GM9AuGx6QeCamjrtDs7YX9qfLT2ANJdIwXCO
XLYv73po0k3VTM9D7iSBQwsclBHzlhIUemmGItWXmkY52ybi/KyQpOkjWXJSr6Cd00y3hGSXgZU8
PupE+fBqrR3kJLzdvpD6Cqi/kb8A3lHIZ39b1EnH2ZvY9u8Xt4NYTSaf3TgaYXhAH3YLkBM8EpRV
VUU3VN7we/Ejtlf8679NhpjFzrNy9lhhLQAc4F+1yjdxy3OfIooy8UtrD7mbf4/J9PjOq1KnzqXL
TX9glXoogygn/z+6iLNTPh/9lWuoaWtMUkNKBUxUoXOzI/k0vfErdRjwyiBL5ryRW/cYIlUUXgl4
WRDP8rLavNBfez2DzF0qtyR/UJUcFUMfGn0amDKfMCzAYrJlP58zk9kz4oobk6WXdVNxq+dYYJNH
j+CeS7Bw4qVJVY3Kx9JFAi/ye6SRlyhAUx/o2MK4HDeK6linzvkigyjMpsn4eupSCXtc5sUl+7eQ
3ehMFXVmhbukOFXu9Tl8Nw668t7znUsatF3X9pJ0hWNONf7qXqZ7v7LfX9Jp3IvYFfGmb7PgZK0g
/h43884VcRArx0+BOxBAki7AlFe04EMuOSGnVkplbT/orCX4rE3Fo51DY/ssRc2Xq/wl5FUOFawc
Yt6s0qy1V8+SY8VdttIcFPMDYrlD1bmvuN8ZVMymY6nRrIB59Xh0my+n013ILxii6lTwRdwL8CHh
Gw6HnlbE/LSxR689B1u7UZpROU+xPdgqPsUIYwHHqNYvtCQG1rjNYg5dZT3q53Tc2y0+eYm60Nc9
Z/h+fSnoj8NLTDht3bvA0TvCdiDVwuM4r2r6iuvazEum+pZtRSc/Yn/YCKH/3WFqx/7tDrlcjLTQ
pxfTQ9cAfHQT6IvX0YV+MFXK8snP0vZgM4hbm2/p9Z/AKatpiCNnNiAR/4B1TgwuKydcF+ioMneG
85vW0hBs3hmH8v0htdv0v8Mzu1Dgqol+TSW1LT72x4AwTvhLv0hypS/NNv1m0qAwDQpLl25un1aT
JUh1Ql7cH5DVwXKQFxaTaFymYpy1TZCydhM79tu4O1bK3A1oX283EXZLyoWSbS3bNlfkQHa8Vaa7
a6dZCTdZChriQCUyxWz44LqV9LmEoNEP6CuNlysXRe6Kl4KiPx+ZyBRiSynkMqy/S7awD5+xc3sF
gfswEL324cXizj0oZ8tR8Gc1BomY8FnjvkkI3vmH+COpgkMmbwYGHZYFyqXKoh67vFi4WpbUms6F
OxrfVMnk3aflVpOFpVrBKP2nRqHn6cAH8R1/PT1ZBFfCxRFpREjjDzM6uxmvo4WevkeeJCZG/eAU
2t+GXeFbKCJNnG5hRRCW9uRhq8cZoHAx9SnDxrmz13sUprpd84xbcQRgnw91WvBLsRBx/icx2dsV
z4PLBg25yG45c1k0MExyEjUba+adw1iukOB/5rlgfGPHYP4RwpaJF0QUG7o3bi4cyGFYwnvL7lNa
s9wTx6BvGpMjZz58tbdIbLKSsPePiWcosDhV7VH0DxOPmImuT9u4QkboGFHdYztp8GHR7CJgMrCm
yfv118WptRJTkSF2iWK8/BzCYMpXhJVBLMaa2CkEh6oJfN6h8wP5C0xKhMARoZNek9dMyHqrmrhB
a1QAAFZzlJcc7CtXNko2yqgTtFRZCCiDcDkv64lwFJr5OoxyY0L/L/rHNypaXTDbW9PIe+8DdMj4
zsR5eVoDRq1HHoj7FNb76Gk4X6P6SiWpSew91Gf4zhIT6whHhNibr9weWMZX6UDHP7UgnLsr21jO
sPle6I7gG+psNUUWsQKWTGxEh8CT0by89N0ZfxJwJP2UPYa9GYRRlC/rYlSQ6G93DqCzrO74WrWs
3qG5NsUiPg2mwLL4Xnx+IajSg7kBl2Iu4+s3RhadbvE0TZX8b5ju1adivnBrza4Z1aD9SjN4Be7N
8Rl/icuRtkHjmtQk6nu3OTJ1igeOSUtMJI1reFuW50kVoLFzL8JviF9aNCEBuNSC7yaN5Ai3S/Qe
450TWdjsB3CbCaC3FkmDrRdD0xKPkss2mMx6GFReNksJePw+TxhOSZPd8CCLBeLXDBiOkulTgzFw
/FOQnhCVhWzssk/GSd2FUI+bSQJGhfR7EsAQqHXQPSo3IKR2RWk2WukfUK7LrqDp0KLNCNH/zmha
iIkxP0QIqt3Vdo7ttxpwq2l+PAaYpjd1g4z3apMruE3e9ice8yi7MizRlLa+3F8MfdenQik0IeAl
3sqoxv0haQbadNnR0WH8J1PYQ2TOCq96pFtoqVVcWQa8O/LLb0kf5b9JQHQ7VaRyeJBM01kqkxnx
yvcsgplchOdYyZQIUV5267zkSC02sknnSn3dkUMI8ciFWlwb1Y2PZymC9LouykmVui+JYRiKtFN3
B1toX/DKQtvZEJ63iu/pIyCFb2uNFf5EmdQgKEO2ztBPAF2g29xA4K11RhL0l1sOzbIH0yeh4CZ9
9FNIBBEUOW+Sv5XZ05TGZBFyJik1xda3i3tYxSNEKTz7P7NrMJytlOolN6M2uFt3KpkPKkDeRIet
uWkOtnOd9KoG4mD8cQPJgDos2wHP2G6AbxWxHmCQBuM9Ib4P5n4ypDyfhHonwPz36dlTswZwQigQ
L0eaFRMkY4Mi5PT2aqWQHPd62ilC9eT1UQnzjFpjqO0SyDUe8zfQC8297utNtGobeEzOWcCEl8aK
lUVkgJrEjRp1DtJ98hNX7Wl8byucZa/xxl8OT0+Nk+5fEXPvi6DohV7GBMEUqZSkgUYjrnFCykqI
TYOkd4tCXWEUJFckDxchYYZewQh0fDti2oRvOBRFBfCVKHEryjPqrXx5p4nvAlBvQb/pn6HaoPqM
xAnYaMM63FD4LkmIunu7L6GBMZWxeB8UjswZmuH0zJ7fG3NKvZRH32dQEaGVU+lF9Qth7p3k+cH0
j6iOtlHDuzE1XKUTTGmD1StXQkN4TVyu7+XR5MNoLrPxSqAeirAIz/gCqpH8iJj9TrNo1B31NKOB
W1AmynORcgfUEKPYU5kLUTJYyXXlotDF4cO5zTvehhsNkrWdfbK7ca0a5Xia1oAVUaxJVDnF/pOH
Q0bEzH6ufqgDRpXGhUVcN9q1M2vfzFfqoLNJJ5LTAd74w1oMcArfIb7JaGTLpIzdss1UZZ9RAlaL
mwob8OWnmc+ptdPAaeEw4X1qCCdwevdm+oqj1oLimT9A6lM9l65cqVCGu15aOlmN9Q9qfP6+/3jK
PhgLjbOVx9uPq4MEDNjrXij+3/GYSJGsuggBIvFTCsFYIcxIsZHSQ5VohuqPDlg0zgoF5COB1wjS
8BdjP16u3qmzMxIUuzS8sPPH3uhT4Dw4mFGUp3c3xKOmCCieIQV/emAB1CmD4fARgY5j0GLE12kU
U83nDWB+a19SHOBlC20Kc1qGhjqUyMXZpIWTgEzpJkJG9I1abpJmCbYp/dpKQHINYu5KaVLrZefP
S1KAJUF5fSjgMJiWMik/NyqbrmDhZ78a77wLQbRJjiz08emT9NClSqF1JtvH92ZIWIE9A7uFNdWo
DwDvUtUBb9kBN7kAXOQFbHT0mxkqw+TmRN8Hv+LDPjmWesHINI+1ThwMUSj6DOEFKoJPoSmUZX0B
gKm27ntLWYuIaSZ7YOOoio1ifh/ZwionoubDQFELmDI/97cAp71JgAQWlhDZEVXd9JuPOVlJGDf5
RqpALwCxAgA+Q6sxvQK8xpvaSDvyofvaufI9DZynSYLguq0aq2B7Ac2NRsTWIKO4p+aKSeHgKJyF
XjZu172hHw2HNOYThuFO4AdFVDSvbsFsQ+g3rfst4ZUPxpla7mU6rApNZ7+O/RK24acux+KCBmuv
ptOAk6r296OjH+Wb26XODcqw/+3wLJWzV/kKvRih33lV9OPR7epNLVcSzXiDUYlXZzDbt//IZrQ5
MHM3yEpDCAi++y9aE0Y70NHJHMG2k++wB2Rnub4RrpTLUi4YkK7YX81mfA+Q//YnYbYsAm0kKU8Z
BaISDieiNDNL2wYtKD+WkhRi0AJIObZtWUioT6HfOIXPs6bHifMZ/gszX32d7NMBIQdnfr0F8ZXt
Y3iplhUw2XG64H4QVZSSsNKdcwvapm/JwZkWbgRoAzMV3PpP9Bm1jIzksWj7GLZCAkSIkNLFpPNB
Xiwz6Yxu7uvrjB0/uO5RtJEbf5he0ZqA9jd8D0WcLngiiOTiTKB84BsZDa8KIq3a5W62zX4mFZOH
PdOpHeu+av599xYXpeiVhEQWF9RO04MlhFDsU99KDeclfgS/MERjx/uqASvgGXoPFOnG+7uowmPe
qEC4QDpDMSRKHBkuQ1nEsgrEjnXcGI4jTcZkm4JsIgQzblo3MLgDtdRifDvLvGb+NJFuYvERUL+9
5OhDKTiNG95wQ8C8wUHvX6fdMll1EZuEXQUEsOjDO/UlcuH2PAc94LxJ3W7IXQ73RI43wp4aJ3k2
o5pAu9xeCPQ/eOApqWgJeTjnQMZ9Ij90uDfuhzeeP+0KzRkruqMBF8TgOiXiCiYNfEqRxStnBW8Q
TCj+Kp73ehTtipLN11kpPlzfSstVNUfuTPILX8OiWfnbTpETclVA5S2WKMhYdAyIz2WDSnroWr31
cFKOOU2u+Yt9rge4fz9vdYBzXgKxWMx5w1byogUSzcPgQPCf36vKvHbLQJg4svZtX6zHquACNGsz
d0aQfaCzqbdqH+P/30nVQt/j92D1EcMfByZepVFcORE8fg1ty2x1mDVb4fk7xPE7TOGn7BQt7jEC
v1wVUrQ9oajKhuURRigZeUn5OCgFkg7w3ooAZ38A0uxaYY0zVIgfrzofIdjq7zGuiJShXp8v4u4L
TCQ8KWKp41KSAlSf4RIkn3dNsXI873J/OBFciDrbUSpdN7SRBFQgM6ePG7XYJzfPa/lD5TQb72h2
JpZ47LeDJXWPDx1spL7QxIGuLLEUW398QuR232MACWAEaXhaQMFaxwC9ca5Yga+UjvKQ1rIfvCdl
rQx8DROy1w6vawqCUuT9GLTUNcRn8xvlCQJ0EqtMIPSX3yqlOdwuc6X35Aq9Ja1xlOLR/FSSOMrX
KTr5YdvblbSWXOAuXV7pcUIn9qDO4XCpSzk2EvDDcTWP81C0B065OJmaicy+eufbzzL+Z2S35T0U
VtFEA1Mx+T9v4n6fHRcb81l+wXDiPRKDiL/l9KVwG3dq5AoLkw9vLqtvtTqdaohZWSVQmkXYJiiZ
Z4vpiKx3/f+MvOjxV+jocOP8JyceUd2HULW5TeepAjXh+wVmnu36HVEiRko0oUvV7Twnc7bTklBI
mmSUIwqmEVSldtxaWx6Goi6SIwKa/7pXqw3VWBqqEG027Q+KDRB2ER/zJFEYSw37oNjK1MiQA3wp
rs9xd7tYcKRHRCESfE+M/Uy0VwIuigi4oVtbFWXnZ+PZlqIkX2HlljlTHSt8ToaYaN7dSn6INpxe
K3PaDcz1vGxNm+bJr8GEr/6UEew7bS8/6t4ZUKrKHAmcLkK3dZ+/LDZjh358rMj32Y8sFzElW8R2
z8j0hOfHewtWegLF8ahx0MrDwQHhoJ5q9MRRYom/N7+9MXoM6Swxlvv9NOjDkB6ll4dipcW6oJlA
zeaRMyc+NfDMaFm4HDWn5GQqFvFjQRuWNP+dWf+pxUKvpBiPJJOqogdHskvbDFVzWLU16YGJtCAy
HHfW6r71kkXmmcWZiOgw5290zwusHUip5nq1jm5sFdoNBzCLhvhZlYh0W480b3UjjWqrjnyOMf08
i+tCmDJQlp5UmV+0Num9/iRPVqSCW26xuGo2KQN68wJ14JqwgoGTroJM6p/8hRCw8ZeN3srqxs80
dYHgqbttRrEOQV0/Jy75zMTkcajdGmd9KgPmnZCmJBxW8TtRENs20e7L0xp52NV1I+TUmuLFB8dx
esRs9d3z6ev4K+gUFcTI0Xaf2qowGuvlG3xB4YfaCSsMQ45/7axsTBhz23bHhKQBjxIYP/MyCzVZ
xJc2T9CKe4fhF0e3LTrivUfxTWVS7h25cxjCJFAAdL19HO03M45Zx/mg9z3lSCf8fMqFILOqfu+5
vCefWqv8SEcGi+BvI8HY082+IQduuiG7afwU47Yzg/ex9HOoxhn2LCKRAJdMtJckbHThSICJTAaX
NfDgEnPuHVc4u7u+OqeWgdafikLYBssoDVJIuGoSdqHxJtQ4EaK07wnqZh13+ten3J2EBFNXXsl8
mjwnEXICQGBDqkdCufrMKw6/iAaXML1pp7P+LK4GXIHYRh0CmAD9c6kSC+NVyPwoX0p0O+Oq4gVF
fpVHAD2uQXvd5UKVyxx2DvJewq3Eeqp9MAL60IrpgFGTHexA9t/uP8YXsBj1yoWByE0p6uJEEHgS
bjf45XNGmw7GYduKJHfnjBaExoEpTAlW+W5xBgdEZuHu53Ld8UkzyLSIxWTEIUqqFaS571jvB7BY
csu/fbs+/gwdq7jb4HJBzvVBILKKYDD0/Hy9yUmJDtw6FN2KjAn1Req1/+mtQDVuAcTvWUVj/KH+
hM68/9sdLvnC5rCNYCMgaz5XjuVABQzWniJdU1XaM1aBuGK/OhZjiXZX0PTwVyyFlutbeeqEbhEg
8Zxk3EU9E1dU2PEsL8D+cXAPyY7Tk9qmC1d2ELhxRZweDCVitL7fAzg/AYzIachgyjLaiDpMgQMx
VWneuXXDxdBlTnrWvWnWsAw9bnYY3Ckl7CU1q1imdFyB0pdORKe5lqKWpC3N9v5ZLmvDyO8qPxcH
1d/LSZKrAy71fKOIlzpfvqJ9/JRNj94jrQo18YraDe1MxYEICm46Fs72Kc0+t+aE4NIOh1QJmrI2
hoq79394NAYOTUlCMMnZXrst/3v20XUv+mxr5CE1ZCSeQjPE6+XYHEbmVBsz4eK2PBemFZNURMkx
MG4y/xf1JbMysGkIvXbnVXycGczknRuUss0TmDN4tmdm0pOj49w3tSbev2P/nJEFsHHshHSj1KMH
tfbSPG7x6fge4CxUb9zVQzb+vklWxjNJpfjWSCJz/gz5moztcZ2R8kT9MngsjaV3kACeOTP4WRdg
w1vN1OPdSm5GfvmFNmkH2gXU844sca+GNd76sYaeSTHogttM3W5Q8pLU1JvN5bCbuByeKD2qi2xz
Cvz5qOW+qcSuBD9t/1k5+O4Rvd8nEoR3spZ80EPl6hdxFIMQ8cqUfFihquDLrHvuDAGoyrE3rQau
YA7KIxRmFKJ37miiKyD9hN67dwUrqHjQJ4CevkBTLLzagoteaMO4XB1ZWjwi9QtLDQG4Aakq86Xf
zK4YZd6MFhgUu76pVxNibjLwW9LyTLJdvr8iU/DnHe8lggjLdtjxvSyv24ruNYFuOB53ESwrIlrM
BJcG0JaRInUmawPUkdSrWPd+jbLFnO1Cid82hrqTg0WAXoUep/+n4lEduR0YPv6lCgOHNPcwy8zG
0v9WCoAuEO0j41zzFgZXRjPt4WEQ+2z2WBZPphZoEJoMi1DgpmSnNBrbVMtV5FBomwq2f3ERQO36
MjvwOmbzAaLz6Iqwvn9lCvRssdEKv496LXa8Vs/gplNfvYqwWALClHeklaDPTOh3C4tr5JKPT87J
VW0lJ5caKzua6OVjSl62WZ7DxlRv22TXsPI3Nmno79QYziA0JlCeoNjwZ1+H1euSbtp+aiELqQ+G
UYooeAld2jyHSnTBg6mRo2hKhmaTJ9cTXxkOgo7BPpuckTuZOGfoFQu7nM+uW5e0o1i09IcMAzcw
88TFPpgLjQabfY3Tb+HHJBw6tJWm5R5Mvl2K7QXiNoEtusPdWeuuAXcLGq743okh5bPuP3eu60Py
Kq2KvGf0KymIf+hZXJVey9sX41Fd5DXVoNOLHk8TnYX4kkwjdcQRflFHUwI7a3EHQgvu5dfV5Mie
fqwBx2BQAfThnrZLdo74U4kTiw6OAtU+ygn3sxZb1A6tD/X9ymn1BViQpkQMVepYuHv3W9cTMpdk
LCsZ10t191MhFUyWFRPrpevj90pBeiEt5bFQ6i2QlI4Zxqw/7B8rYvAgSsYpqqgW0wdNM4urz7sU
Qq3FfSDJ8ymgjyzhX04wg+g3zAVbpwuWuPmzKbhShu4YLrDflwQF8i4DjNIUl9UcbuhLJ7VWeG0w
IGVM9OnUJJMHGuj14QIDRZMCTrazfrOSbrt5pq/TH+rzw3TJ9dpxXoaebgeeB3nTptJsyc3Jy02W
HcmklkGbWDDovgNqJbrYYNLZI5/KEOqGbdYo6Yc5rgj9cOEnG09RFhaenk9mSp6X74LWSxO1o+IK
TgCDP+kiQQ2M0RkhtvXqndJ0+lxa+SDtEqNByyTP2L7y42bPWhk+xXbNQsRq+5jrphfo1zCBDkNf
rttURX1uGwDq1vF+0GpH0I6cna7mN9rocgeZAim142IvvWusM3BWq4Y7ezjmcEY55VMFdp6XF7C8
HwcC4ARe+RPPFJppwqC/FEgtqTV7W8n80NSwa103lg52T6h/j5jZMdGYIJq7AG0GyemLaNJ6jjRc
om36VJVbh720b77cCxeR8/W1JvQ8eD7CvMHLRv4lS51E0kr6qot5pi2XxScr17dDVA+mX7ls89jA
CfEldrtGCsVHhCcPZQyhAIYxkmSLBTtzULE1gkQCHXf9L3+bvcqnYJHixa0zcVHTieiSF6TRpq9A
DWHn+Rhcf/UhFub1SuBthfDEuRUSOt5rbRiXiTi0BjQsGI7nGYEpUiyI1/OF2lm9O0uH3vcTdl2d
MJjErKVi2jEzqZk/dEQMD6sr7ODa7e8oaPR+HIQquC5U4+okvLcF7asx0GVk0boQolKHjWcQbFh2
vJ2rXy9O0Yuy7NBemehoBYN6LFzX4PbKjNith8own5f6XtjaimepJq22RClfZ8D/DlDnPB5Rvl3r
vfeC+LR8fo2DsX5xaVLm9PArdHFUuIUQI0++bWvp6iEeauMALvZVE3IX9eM/zdfbqPyaU/1PbnyS
+X7GGe2bb2DHjYWCTxwtmrfdhbQe41lxs4upPRiEAR+55fQyLDJijsiZm3bvv0y5cufZd+JGSvlv
X1GjAfsl8l78W61yOkTIsNFSdiFyWgP3d2Mj66kK520an+b48J2Nb4qKyqw+1cHHxVl0aSnAktTd
n1dRe5FOUJb/Fa+3PxVUqKFnYqiJ29JL1aZQfaqVG8KFNkTvcLjF3lktWsH++L1DvRsEtzUpYfke
vU6CUBQNo/jIJ4Dyo8g6bfwUsr+WiWRbS5OzVCDHFYohGd5MUM5EUXjBuC0lCSJN9kQAsRX2sud5
UIcKQXevhrDkwh3ijZKrlBAvJ+tjXTYoUCOPmzQJk92a/ud3tgdQbD4N8nPHF9WW1Ys6KzS9pdyF
Ayne+fsfAdv9Phnl7i7gFEAW94SzPE1xNdCjvn9Uz5Mjzv0g0HwxT6YBzdVxK7+Kf0nd8neeQwHQ
RTN2OJ2CZIHHpOWMElZPLaMsTHlSAbMl6Iaju0cGj7SxbN7pMqkq86gq0qwXclN+PtiwdRcITXZm
lELFfiEn4JSHG7/ZdaYw1le6evtc1v2hlDDG0gImCCAfN0VYLkM99A5x1FrsPm8+Udg4m8EeuVlF
kb5T3L8qbiN+l/Js6Owpy71K7fVBl7nqezV/c5nJMoIxd99WbOyMy+Sfqk73t3F0M/6aLH2fUj9h
M/sVaEeVMbHJzmtE/gB2es1FTAGa6BqX4affrF8jOEYPreUAvB7ZAUfgJTtpQrlx1UxTkiCZzpYC
iB7DHXUArdSdyTwCQgqXkTNVcSF8+Pdc2mg6iUOsRQ+vyUCsAsqHeFKE95z/JY5+5UQoIOlnvPOj
czTpsVmTCbVV0E+2PNBmXw+LkXI49TOCSXgcvv0MXykKk4qk5R5azOD7Ui+ini4vtpHiG1LnlnyL
ECruYbl040onokbuk+E3RHlDbXOLdnD/C0iR2NE5AkJu9kFzj2y2CeMBs/TStdO1jXFhLXt7Q5Sw
5uFb+pQ2FbGY+3ChWikV+1gRHCOsnhCBLPsppPpDRF/jF8RXD44umpcp8kJpJDAzrKtG/pnCRauq
peX5axmaFLrSn53fJ6HWTbUjG7YTYzkaFXJuBQbovkzyvT7pZBKRaelrmvTd9aKqE0x6njpAgaEA
aOQjGGbKde5SHgOAe7oFQcOLx65+LToUoogH6tp3ER5NTwCmdwFNk/VZTDqk5IFc9tvotGf7Y1nI
OH02ng6b2JSYJ5FtcAVsDhvNKq3Jx4++c0HYZdo9dSeZUTuLfizHWhJFZ3FObVFxQFuccS7htpNw
b/3cMVC1xRTHEeFGLEibhRrLeA8Mw6yCcIKio+7KKqNuobjiDsET+hrlJlB5K78aMyPgWAaqviYs
lI96tu/zCDcf9jqN+r7ObnKKWWXvrHlrdGyvJ0X/N3oHq0WFQfUIxUOi518vUA622xbiGBczarWd
1M13LKVata7fgdmcCEGlzg8WXsX0jFjg77t2iRF1Ngpct0OegRonbJqQyWn2UK4LWjGOJ2Igov6Z
HVRz9gEwm4iP0x2p3acj03o+n+JJy1kilXOWQJkIqLzSE647k/ErQ87bG7sycKo61odOP/v04ES2
gp/qwD+IroPe0pD1UQv4Wh+9Y2SZowNJc/kJA0a7Wf/Z58R31D0uPCe3/O3av+V6TOWmOAA+NgFW
z4a/JgEW7pmTU2UzwdwQLe3IpdHEv8IOMdzgRhuvB90rKSIE7ogYBAIkiF2vgCeff3GULOHPRqQx
sS1wv7R5/4U5NNpIz0q7LDOZ136nKe6uYiqDHuRccA3QcnyBM7ff5YBzJKI3xbhzuEtIgoZ1PdFZ
dEOZ+pJC35cnZ5MDoXCpEffTkJMUXPfGh+t/XKAQ43BjQwu4cMZnTb8FJjseanEx3iNK8x8vN8Ml
MqJGeYGEFsK31nKneiT9tNZH9DPFjzVy/g1LvC0ZZ9qgdF9DdPrZRGy3V0O862Ko0Fc1PYWYk+go
XfMez+8nIaFilojhs9Wogn9xR1XLeUeA4TKUOp2t05k99KSGDA5edyfgZfMTfS5QkG5AoydCDnfr
blnrYDtTt4TvQXY4BlLrYJTLiyBa0PnDB28zWXMFEATlVt2zCGV2ru+uCKkhxpKVaygHICxJmNhk
R+PPl+LYdzwapEyzCtLQNiNQhN+NArJdV4RxRtuxrwfES0QKLNIRLhicwINVD7A9x9Bx7ruCUhjX
NO7zWXh/soJd0PMkP4n6Mw3VY2JK04KA5B2srAKdFXNxEJ9jRsuNWaaEpdqnENSFejI3IkpAWzEp
PUanuot7i+qwBa1N8/PDj9VijV7QTLKom7m7ZPcu0KkGv7OWAjbzYFxeq9+XTXgL16/7xyzwcd+J
jJg46elDxCkRtTI/PECesrPpm247vvEjN2ZK468H1AOvKZhRO7uV+Q5GkVbN0FO1h4SmQojKJPhS
HBYgQtEJfp1dLeDHbGuhI6SagVH8ir3lz4NKKURdB8Pmzp8S9UaeZrcBMcUyuMCONwSMt45rGpHU
7N+wKhSZUSiUuujOZ9qqt6WJ6xWgC5vo/xohahUfGDlqeBBQYgIyNlFrpt99HXlRgpw/PI23Jyml
50KJs0yrm4ML8jLddCLFy7pGAUGTQXxnu6Kb4hg+qSq7taaPwOo+HM/Cogb38N47SpiPfIFA+ocv
5306/niNa0vRcaPvroPdOVgh7A9TgOCPTHcyiB3hnAv6CI/oxpBNj8W9l2PLM/8rn/MoRbSkH20/
P2fcEDu/7vn6Xso3I+ZaDBdcD3n544WKrNAqI5k5W/qb2in1xbVmaNu/mb/c6InTHaq/LAIV7mPL
WSwL0ZhoGyswHJLPhEaX/5HixNDqUmgPoblb22u9JNctUxTI0NBwfFC9mTaXniVurGNObm2qSVvJ
Micp/xIFn3HqImnpB1e1ZJ+NgkvVRzyVxEq9ggL2di774f1wEpa5m7fHqrjQj2c7vwNLUVJ65oXi
IA4XTMRBgSIF1vmGZro5vZTumhaoAkJjiyxCjjSO+AW37YF0LjmLXRygGwuixW1BwvoLZBF6qmEL
o0aRT1+y9FS5JxONt5mUPH79u4a7mlDfFEscoVJpPewnVXaSymE7jfeEoc5lkxe2wDviYrqCy3nx
kjxkqvyE573AfvizVYgXMvjAN5bg8uLUNT6C7JtnNv547utgTRVyC+Mw7b0IFSFvcbI2OBZe9m1M
3FCvRQLjsms4Cii71TFGWSmVnbM+uW4Dr1q6HNw93nJFIXJxSHQe+wnGcRjgglfkzL2+o9YntLo0
YUhkXOyuOW7TjT5w5TW3KbxJIKZnVDhITXRtmjjm+/BDwje8b3wCFhAt4GA1iuEtAsOp2l7Lmomp
i6A+E4tMnThRFoc7YFv8jOCNHJt38dGSmhuvRESxE6mHz8iv+4U8FveB839fLkkpeYxBz/zmt5qM
fQqcoBwaL9l5CtjioZ6gPjT/3OpEaXN70r75X8062TprzZMUm7cogxp1RDCXxbe36HYZnhHGl3a9
5Kxavebx5KnOg4kAgTyjYu59s1reZe3Y/bU7mJbSU/HR0ZRkT8tTh+UQsdaCpey4+K6dk+zDpWqN
V/mMNcbOa/rJlIdXp1AIw6MyuVvqnn7gfjoO1aSndf3giJEO9OUfug3sX2iUlDgi7jJ7lHVn1JIu
jmaYARPpEFVb5JusmL1lsnXRB9ypy7UjvYgwCrMAl/T0HoEseVLPBgM++/A5y6/adZAT1wd2IC1g
EhLNnxqVmBuSnPvOrRnUh3vkFOOdQo881W7HclWyvBrUaC07ivEiMN07b6WtTct5IjheorXCz0CT
CqEkil7dfCT3bBF/xPpZjB9u+vSrVY68UuMBh8eOCFqFx0wuEm+EM6TM2kZbbIb4mVOncno4zCcz
e617pHtaAvC3lqrGyrtvhDAueakT2QUbAXAH4jM3lKPRqwsZW90A01SKJ+NQvLvA6jG57r7l1t3b
v6yQMz87NmA3Vak6RGSFW3N9W7EIir9YrcE0RSFQquGhHDVB80ItUt0GBsHexn9YPo4vS8IawDAH
ALuVOgf9CAEd0t40SNXv71+8uagnaYoIMV79oXpKt+hi59o3smwZlQj4nM9oP1XTf4SMlZb2DeKV
i1r4xoKEKcLKhqA++q/ysJ7uxAEXX6Sj0gUVJ36BqBNs9O4AD6Yrn+BRsUBdtT9jgmv83AJvOr9H
1EdygSXF76c+oML1/p9YX5CS8bEnu7BnfW+J1kMdzRT1rCefT6Riud2PNuWDbYbCkOInv0qLPPNt
MwP+tLS/9zil50U2dSE6E2GW91B+eQDT0M+kMBjcL85E0uY2ddmSaEuVG7eMfWFQ2AvrvelGo3yF
zXNPTjJo8R2h5p4gvjldQ2PZbfPtKt6mop/mD90M5UmzmBfZsiAJPvTCWakKK1kZoz+KMpQFr8vj
njwTIu8I+Fh/Xwp39T7/4+ShPYb/N45afN3wFqVTWcB7C3MFXlvyyYiMXCTrvP+ARR0DHHndcwym
Rl9hMGI+TqKukWCSHDQLZdJie1VHh4uTpvUnaTqGsbC2Wjw19w5sFztRPRL1A+pdvM4e+Xyqu5U2
XXtdYYCcYeiNIFVeEom4Gza0gunchNu+fsDDwSQH5vdTFBI8TFRfzIqkUFLpEK+dlMdj1+uLPo4v
nUvnh4o/jwou3RGI30qpXoGaTJAfHiOSKdQCK5DdHooPmZG2F4HOFWajc7VCVrIe7QENMQlTvhKW
psRnDSvjqo0prA0milU4kkIKb7LTjaRGylquuANT1FUdPn3s6yLRbS1At7VjlquFUnWg3j2Sj0jh
1lG3gd253/GgioWPybEG2c9PXjhOcScffL1uIggyZcf+PeXdPQcwTM4U2k0x4cyQ254LGD8wC5Vk
UxdEZjf6hhRovWRJVC9wTqveUOyl+wN6DcRFbFbdhaGHqms4WBXQrWTOuSNEsAQLS7VcUHBg1O0F
v5J+kp8FKUl5HYRlD43p4WEAMe7NMgY6D00ELhhba1L2W1Q631NfQDTLIcI4HAUMOR2V2VZass5x
NdmaOhlkAeXw11mAIpqW+a7ePowwnejb+MDaVSmLVNNF/KasgriQJcR+1klV7ktrA5B+kOYbsb87
gwrKPBbNQ2Uu5o8NZJ76reREnF4T+BzeWl9H/js5lck35u68h6Zlce7LW/bBnZAUS3dtsRM2tCx2
KSp37DtTJtME/IlBBSVLzAoGNuM811QwXr9aoxnBrgBC3PW7nVJWsSnMqjq63r/gOMypySO47XVv
f3ugFbb7vjLHl543cydxwhz1KYQBYJr/1DqBlJZgelkOVZxocCCozDJTiDLqAIx6+FCkPNVbIK9u
agSSSSW5gpdD+cZPouY8Lo6NNavKw0n9mhtbWJWeUm5gK9muvC57fq0EdBbk9le7YstkzABsjnGf
DF+F5KQvbaARJtGW+OoDDHxHW4wuE9xpB6XhQI4QVbu+mcEYm+UUfyq1i0emf8eyHcgNEVjMvheS
wBsm819uZcdSqTXTwgfm0EJ4aXfoFJuEnN4tPC74A/JXhfF3v1qn3nqUhlc2hDabF5GvrI/PjqUl
8fWG2YoUdR5KqXELdpsJG1rwHwH2e6WCBIRl1KDr6+FWCDLpEv8ywvpZ7mwQcn9Ib7AWhObIjiPC
rwlQfp/nMIdbVXO8hqSQkJ5kXwtvf7vclyGLgAeEG6B2DqU6jNeLI9McEwYW10/HeyxKkNt310Wb
K77JB0Zzun7LcUQ3cArB3+xsFPvg7/ZoNNi2KSKXteJAZgjTmUZg5gFN/v0m3pRqX+tbbq1INhVe
4//Ce/krmhPv3N8HUVgdqMct7inCnEW1VujPL6wj3GFsrWsxfnztZwnC7vwq838uwCtoIF5WP++2
9jstBY5PNtJd1IzYWTbtDy4DBWfBTRaoKOHrcspkyL48YohM1PR5XznB8tUpG8ZOabWgAb2cb63m
PNJfbXXWcEvx5NWtCLRl3coDsnGp0or17la2hv5zCaH1YjISWMzUEn7jOSRQzXAbrUrJe9cQrbjX
0SXxtWFnW9bcQrxyjQNKpnOdRs5dggRUL0z/lZdpAGIcNPJ4p6PtNw0VX64hYrBjP0MBVNbZRb4C
2282LCx0Zb/F6BT4jwl11YWAWPuO2mNytor4GIemuLbK5ayWJQNu0xJH2fY3w5s0GLVaQGNiEO9W
3BIpqdq8l/WIg1elcJPmYxh1q4c5yaV959fmpyH8rA9gvaKHhJCxB6FS++q9RvG8Fe3THGU4muEB
l0x4BGJzmnsJmIoLQqigjSX0wjNbT+OKfdlc3lfRAqm/gKgqhdplkBXAv+lYy4jo3svnkBFudBkY
8VcPaPpvZpMfqPC5BNDf+T9SFquqtHxvPWs75wdspbpKgU+fUkXpm9mv2Gjtu9a6SRMcjCX95haq
w8cSgrhj4aAN5lE9l1yFtiY+IWhxmEtw5CytwMkpUeYVYrXBwbF4/fcB68zs/iisqXzCnxbpXmU9
VWtKc0xkJIQv4cAp6jgoGjRKaldM/SkccAEKjQlcaE1NRhtiBbsj0IozXmQAzKAbqpDRq/GLkrIR
FP1f1n+C9E5jnzIWs9xbJm4Rm8iTf5gB0zJb3GjSpx89pRJDO/S/Hix1usx6BGDlW1PiJ2BZd+2Z
ohFCRpT9s+mfgYY0cK6bPj9e9TYgfdkRpXN6ngD6Ucb/NXkyrMSI7oYeXV/+KV3ViV2u3bFFAS7R
4dT3BbeyC91Hdi6DNnB+jgYcH9y2n5XY9NQTIe3FQDv29MjdMR90PlyNP9LbqzhfTeUfMMw5Mb7m
UEF2LgVHxiPfhQFoniO843m2vLzp44weOMGoDexdeoIkbZShqQ3hFriLq9gIJw2BmVN9zUvLjo8Q
vlWNH+i9dkblSKwI5mmkKJP/sEkUS+ooy8D6Oc9PHrei1mKljD8QJj6X2fAKMEjZMPgt3J9SHmcB
XSY8t9v/1O40YTXbjDz8JDUuG78GDvpa2lqEnFIHV/3yvbs5fmG+IvZ6Y+8urQ2sCrCpp7p/RHZx
M49x9I8eL9rY027W9vWIhMBnbH/G6Yu7wyin8MQNCrQHusmM9fLrr/qOr6DuqVmXOYJY+JxXLwlG
RHAJkkICF1kDanppIGKGAqZhZhT6AbmM2oXE9NIBh20nLsMOGQ+31WPHj7LguXQ0vyLevfe+OpcW
iqqZ4rNJOvuq/xgrTgilbo3u0OiJbBGMJ+bfKXGhICNy9dWaN3LGmPO78Z6/OcAGd15sb61lqK08
yqEPowKcRQBFenNPa+dXmkPSG+O8dcXzIPUStwJ1SygRP7iZHT5qx0WkQzMlexz0TtsSTC/VMNU8
kWZqJso1P8EzoPQtUOvdgH/Umfi1UghPZPxE08ai3vJh6QG9FEu8TQm4R18EtthZd3X8uAI7GjDN
SwhpBSKeq+6P51JlTLT5ZwQiQautAtTELmUhvWkJYxPjthVfpkBbUbLM07J2zdsltOAgkwh1zQwy
W4StgPYZQwr55qP7T/gJDGiZK9yovGXKOjry9d3GFpJYpo8kzauQ+thkStwaKKkLMkY3QiHU+7vC
uIoWlN+XgT/eSw3A6PPcXF90PcvTUa9ZMLfaBN7UcL3jL/KEGAkMy+kcLusX7w3rgmum7Bv8XALG
NzXzceWqPvYjTMhwJlgZyqW6vEhHbBs8zjdJ8WXEfoWiOY0c8tgNqfyjm3Dcmx1ut1gN4mRDlyj8
XMfulQftJhpLKtMsDS0hvM2t8g7ZbQ4IqPYaRUzC9WQoJNUrLzh02aQxaWTQU6y6+9CM6iIgZrdc
WF9/Ayq+FoIdW4w8sp1PWkUCl/ruRJe9StR/MaktMBrRp4hlsQLlcSGLxzYN4lxVVeUzxdZPjTMG
QoBajyIbX1ApVUcywW9CT5uDJ+2eUN+M5pdLNaW5yLyslXm5nBEJWr+iug7/LkxAm4jEapaQUbDy
32CQOZG1mUtyjsIxgQwZ5n7XTeDGyytjr1Y1fpSj05aLGvg44f7WXXLxBX5Fo5Fv/2vUNg9VfPeI
7qvkUnX3H+CeGaHrOEGNMHffzkKfaX8HM1dGFnp5hdR7v7tnWd9Y8IO4k7OBT+nP6ErNokOGNuFa
HyNLgdgi8+P0jpTzBzHL9jwoOtcYJ8ayR307QIUpvrjnLYe0t6S1Lipp2BYQex9x6wBn2HUxReoZ
OBMUMy18mm0kr2gPTy3996PY8Se3VnnjQVTnXaNwSEmWb9po42bdGglCjis1w3AvpIigo5wz2MRQ
+gbTD4kfsXqj6wRKR6iCBYDv5y9g1crvyBJAWlgrehgEF8ph2fStO1BZ5XlUTcI7GX2cGBpw6Al2
bk50xsBB0Sb1g4tKoI0lflZDQPNXVQ1xLAMcpuMRwdUx5WgRhJpG011hb2af7ywkmEXXaaYxBKkc
kpAF1Q27E85tnzgoRAZVyrDbOvBf49PXIQiXj3A+WF3WRmySqjUyiF5JfSRuoWSuJIfsaopCWC+A
1HgaEmvvCenT0cV2xpvoXgK+5IXLR/9ygq+0lDrvbZ8csy70Hx8GAAH7G5c3YcvUdWTjABnpLnKd
Xvf+bCXhibWENzU6s8UeEQ//NLnykP5hRlDdZSdF+XjrFSTfXIGU6WUXU4nRKXhMX0YvndW9xMhN
NlwvPwIE/ZLJWaFBF5zUkXL+rIB2HOxYZqef8InY9OUYyfIcSzvqNlepqUYahlqR6mOxitPFE7DZ
PXikXwILP6be6b7+fFu1rj1SJwPpNor4qJrACNG4KIuT3sAs+k1x9iI035MTh2lNDrbfwnZSDfGB
vUCVw37V4yk5ubJeq5UVEC4RBLBBuS+3I+lxkspOJvYzxQNQKGyBCz5b8i2CjI3Y9iqutMwIn38e
EQYFSR/NQf+ZXd/HCN+mBRPjUdSRZCMmg3/bb5hlSJM9GlrhmC2R9uGU9QynnusR8Ha+nBHWvjGF
fnchK3qq2NbfoU/K5bkzfEbhBwZZRTGXIQj+Om+21fyxJSPHzsAzzraxu7Et24rpiPilYUNKoBrW
Jx4qirVEv75dQsxtNXlIM/HwecuUB3iHoOFt+G7uf+gEuCTiY2qXrACVhO4zwZSxLFhnvostYuAm
nqgsue6zHcJfpF4JuNUgbBUFH8wXT1Shfo+0UmjHJJP+pISRn3gzsnqfFCQbes4Mo8rgUjv6iCS+
sAGwSb4K12ek3nHx8DKLhuwzIuEp+f3Yw9iGTHowHIojClZ+lVbxE4WzTDsCGiJIKjQBJYRrch/O
4jQsgwbzN4xh/hYyoxaamnvu1lnb6mP7FIbHXcMfCEthnNxEQddXn4MnB2sx9ba8ZTDD7TKaRMTj
1r1w++eGC865+AUdHxLi3ERkkGpbrVaD1wo3sLM8xWGiA893MM5CcksYXt3LUc6Y1x6I53xBogvd
LyBEt/m0bAEp8UqQOqL6wbOqvyGyH3b3kKP2fjua60/cIaaymKz21GvweKdQ96B9TabcvxnCU1kM
q26uYN/i73Q/RsWrkOsZNsn3etGZBqsVx3mJL/YbMOCO4b5O/7lz3KjpmE2r5uDexhLfFWrriBOH
mKDNbxc1m/fJZjuBT0EmLWZvQVZs0D9RpOwkrDiprBJb2u14GeMteRfBs+j4EDKZYawonlSZ2sbO
t9Hb0JmeLkl01kTPAo4+eoIfwbJCcNGzBScStv74kWfRFHffOH3eHEj58aWnZrxwHNJc2hrjnvsL
+ZpQkia9an2eN96bM5SG3sDjvz/eAEweiab/KMjr1QC/cYYEFvf/RnQPt5qC5LpTB88Hf4KlROEW
PalwCTiPbWj4VAZFy2RDNOfAbz2MBlQOzTT5E5HN2jOMHydDzVXYxB+OMSIfcCdvbrLkChiPcF8F
ptsgg8e346DdyxrAvdJlH9rvly1pNyFlGGZvNWJF5aZjqCHuJTbqlCQLYgrC9gd4RwaV0GIMXEAS
XIvSF6VSGSADOhapTXdlSm0bSNQ9wI05ZqDrtdsTnRnh8490iAxQ9JaYP7tZuRW8wUHsdpZgfgUS
xP6nSMQaz+vk5Z1UCWw3ZQesGFZfmnkpi9Ru9xn0jAj3Nig6bgvwA+JpfTKHg7XuhqZJP/4yToEr
/ZRxM7iN7iV+fIXBXJPXdPoLbZKtiK6rg+i+TpSset7RJlTR5odulgzRlI2NuHOovzPE/cUFg0m/
dE2FHguJJlbIL4IwQmFEX8NTnrSJN7P48kbcuR27QMt1tzAwxqlFsfd4RLx6hNrKPtzgy1Km3POa
E/NdBrBiOQaSaQv6xRTp+8UdlmbbiDn1e3S6ibKP3fBxlcAuwYQqVhbe5bLeyViGttCuK4UU7FgZ
cl5mnQQ3cRyGFbTrue7T8w1fCuQZ2fObOeSklY/PLlMcrh+K3mvISjC+aejLukDkunje5rfrG8nw
f+AhLZbK3crPPFR5JCOJJjyQw2F4faol5nQgdiePzpLOVH9GIrUbJWUCQOhsozqhxXylhzYJPFaJ
EefVTJDxmLjhupid146kcB49MLOIfW9uksiEY+PzJGJqGQPZvFgZrRRtGgf3iN7qyx46tqR58ldf
9Ntb2m533w6c1/iKeEjxJjKE8MbvEqJx1gj/7HMlNpzpSRfre5kEDlI/DWv9NEygIkDXQuRgVEup
tjsdmkhpmPoed60dNGoA+jFE3wPvo8dEAu4pc1PImw2DeKnm0cC7AIC4q6xquTuXk0y1JOXy9/F/
kailX2723FkUgf9JYV12CCu0yBJVHCdYY0ChhUbE9SrDVN/nYIRes6/lC1HXv4qrlDmwk2a2SDfh
GPEb9XQp431ILwuTYhcuCYnsyh+NMehITkOK3MosRsOWow/+A/z7hP4MG9CSvgXfRJGH9itvh0Eh
nCCujRRkymTzpnrmVwJyV3GmZ23/y6Rne2GEXFRWmOqniAP4xKr7Y9f4Cs2iG9s5g+iIu1MgnqGI
rs97RBMPWsJhE7NruXt1ikMNqGDIFDHqNFtcuUrS4kcIMDoqkKXgyLP0fHvcO10uRQhYhkpdUUfB
rcdgvkuYZc5SrCoujy5wH9zk4EX6X5itlZPTeZh2v5KUzO26y6Am4eZSL0SuIqyuRbWLUgsAZtJF
B2f/qUHk3cjivFzh977xQKeE+Hvf73gGjhD50/bOKOA7TqKEkzeAL7uAyo/WcV2Hoz8zCLwYL1zP
mHw/ve+8Mlu26OdFKEq/G0a9p0I254r2N2qRHbGebBtO9BiIAdl/HbjaP9BbQQoMbDU/X2hwElXW
YaWx7ZA/Ym09rd7iPtc7NJ8KeQB+7Xo3prd50NbBAkmyv/PfPQVixSZMnKgBEAGmltktlkycu+zQ
0sxM75oPbbT+OB8XL5fBYqRbu01uvpcLf2CGCJLmCLODT7GRoLn6fOjObPBwBNfPG0yUlb6gSw5C
CFPYOSQQvMS4d0NQAkSTCrZFFmOH3R7IbbfMNVqBUw/nBarUlIOOmZRW8ZLkTG8Q9zpEaPemXoiO
ys/eJGA4lOYvSIC7eUnK7ZhW2TCyR8stPJ5d1LQMEpFDtTU/8ZLi4+y6nLEH+MRXIMvHlMLDe66A
jtCbBinor0SrbI9nkhOjLrlhaClqHbxya+Hl3Bv5FfrX1X/HeHeERq8bzCIfYPimBXUatYd9BOFR
AY/XJGJoSKjfCOm72uRxvU9JK3y5BeeeEHp8HMFAFYJTAeHdrmW/YdnXCH+1dLMdBen63AXwDlBJ
rz5nrS8qsfRg5ZKevi9aXGWIiOgYuUI8AukFpV0MHINEHJrX9+MISKW37Nu819n3Kpec4DAUD4jP
Dn89kBSeLjYTf5fn94xZw60GAIRzMaGAD2FQY/0WVZerV0GBG4ydYWXl77mBd6F0MpU1egDeYdR8
0cXwAgpO1Ma0rpTBirFD1CRK8iUMmgrVrexwgjrXtG6neKZUvxEMq31wC8vOVNgVJkEsq+KFC77K
RP1ujfOoZ/TmvEfa0k4VkvJV+OdSfi4hyGIgMn6LUtgo0H9rtIMNFQsrPGJcpBeqeztR7ApUyNJa
6rsiW8C9JCQd4v7EfbsbTHjPLOxq0WfMmXEOw6zY5vDQexX+BmMY0ZPcwoTnFlU6Ki4PtinTgQfO
dcuclijEC0dflCmPlz/wfKjwDeR+DtTNwXzLLWvcR98CN96M4R8E8anti93ukM8ctFqa/nw55l0d
N6+ezfnsT3a44+pinQxalSp0BE4DASWLPplc6fgZBaGJVx3eeSmddM2jQ6iKzS+hfJ+do18KIbTY
On1NIXdIzNvgZzTT8eqBFmXip3XOyOkalmZbAai3fhTbzXbclTMhcaLdWu9DjqVbFsDRv5lpTUyX
jFw2J6nPbzVtkuy2ATahUkabZZI2/yyXGGIwIeHMBOyVWURrb7RLfkcB6h+L2jX8MX/VLND0Zp0R
dOqTbLR/k/VbMJSQnEFIx6bOlOzYqe99x6BJU5a0M2rypdKTvhaWuaQvaUzRSuatTg5DEND3q2XR
OvD09y7o2yA4Ox1dB3FFoZ6WxNA0OB4+225+RRSpJCENoi0S7tlHqHSgf+1vo8d2i9piBwxYeAZX
MarYX6YdsAb9eHGQxAX+WtyKR2UKe41RG1kL/oraj+FLbv6Z1WJGH07TgWLawww0r85VJpg1n7o3
vfrRjjQqfTkoKSVk46m5B6qHn9q7VaZYIt/6izvU0pvNYa7VQQAoBuVyfNMt7rTJBg0J1s5qM0Ov
uhbvhYcMjs/WIcg8bYrhS44r6ek102CZK/p2c6H0MrwS2+niniAq24hSk6Kl6ExEL4g3soagdYo/
mYPx+K+q8KVs5TwQdyyyBsOWm/pjodAwS3QH9mx7+LOmXni4ZyULMA/Uf1//kFA1Q53hWrr09BpC
uqYOYDPSMll4pZxC8yaQtc337OK5OxZ5SS0+dVHxTXiEicWEhXi+GrC8vtDiP0wH0foHALYug7Ly
rRQCnCUd6GhGRdGTI/rNNPVyt02rAWcS3DtOQV5wp3wC4fxBroHb02mKYn6OckcxNR19acuykkPg
jjLNJcP6prv761w/12OkKpNrJEm6EQjx3mnC6PZQTFMbR7MmcAU9MFZmlivBKnCA7KdF0UC/l39E
RcMtU72KA4IRmRiWAwBBNZynOxnzaI0Kto7UfD+2JhiGuuEZ/PI8NJqzxoGMcY02qg2un3iTSCxB
N/pqaBC5hHvq84VkBO+PRDfPx9MU1XDKtLNPynyp+xjbddGkwDoezwX2+//kObYua8f8QOkF+PTT
AHbeVrte1fuiIdwNSlt5Nk8BoZ1PpDbCXvIEUWMD8QxwVVO1qXw7ESTuL436R0cu+Y5tJZvsscPb
ZyK9oMUYTbb+WkrG4zO6UN/it82F9VqulU5t22S3TyvKaU76tIVB9xXXgUwNZBqey71MQ8tHv5mT
XXqaS9ht+BH5s87mw+VSwDkwQ0YdYMy8WBduwcjcAz0IOzS3AqTByfaHEPWUH3V6jyanTAY+OEyA
xhw/v0jx+PAVrAXhNFoduohMEGymiGQK8ApSeEBF+BfYpsdieu2BgUeSq+T3PlQzUrAEmPBsteoR
9oP1eV8SQoY2LLs9uOldwZta2UdKMlZs7GZIfi3AfG39j/9C8fji7XYcLGQcGWsyHlnx4d4G0HEe
SAP7RJXaPTZyC8Ox8/kpbL/kY/mZ/WNpugDFgHerrUcRcQ4Dvf33VqrWcU2nJDiCngADY8FXAdrk
l+DSQmCGdWDX/q/pdB8QQ4tejx8O3GQVWJcKhwU7pqgLJYscnw8cIHLH6er+zSWCHsHhuzFbUJVK
lJgNmD0HSDzPvaJbRljV9N0DvmdDsBarrwLQKjlwhnzaPEFR3V1ALQJgC4vq50MIRZTfxvC54tEE
G7rDfYMEBxeozuStKn/0lM+pMSi9K+X9jluxsPDwcOwVGSd4OhuPcTINov/jTxlY4ElEHM4KFZl7
Rj6kdUferZmonLFrphvl8gDqWrDN38yCh1Rakko+f59ZKRzRZ6hW4hjZWqCDSe0rsZ17mTmJOhiM
9U1U5J8wApphASADCbh0aeL1I9A3uhgUGtMyERm+Ao8+BAFWwnjeCSMJhE7jCzGM7+chU5Cu34y3
zyCS2jygmPmxYkoHeYYPYhel3ihwfMS+KpnR4YW8rUNMObbQjH1mEcNycpP8NYnaHy48KTY1tyx+
ECb8xhhB//q2dYaKmmk7EEoKr0WpoPp7yWG7v5VamodPLLpfsXU31iBe21wIE4Ec/omsloi6rV7u
K+T9msj+k43oe8SjFSrR27rCB+vEFE28Mlf2I9sGWEfX4+wHbU5E3WKnQPvTmb4S27g02w9LsnOF
g1xwJBVy5ePWlk52vKv131erl1toxgMbxjKTBnjQfK5//tVGKszftzGK9x0CrEPEYc4wSAULWhMz
OV98FGS95TacgjhYlsdUpAQnEpjZwCM0lzlOeRYtzse3qC2xzLWNHgTaes7ovilD3jE6IqhbEdmw
u/2ed+7MivyAzn6J/Gg+pKf3hzyxrcwvdhOmJ6hNsn7IGFDtRX5q5pmsFc+WS3EwsYldYZDByeyr
aBnzsN09l6IM5fcyamSnp6J0ouhWbUpyfx3mKxtdqcOf5CFw2nMXo4thr1TJq0oajZoktJ1DQ1Q8
f/5ssk/LeDJG4v+zXDIx0tRHUUPMZ0x6huNCEg8xmzauTc7jBcyNnpqdHMtpmitzRuZDtNA7QKnY
OEf7CMjdy7jPDmTTStgKzUq7It3npInglSs9A6eD/X0cvxV3YK60rT8/sp3GiK3nt3fOQSbwyds8
o1ICnehorOifq/vArAFxniWEmIO637oByLYXR+ioq5NGkTwvrC3KCWZA34aJEQak25Lhn3hnEHu+
2keTfZxe/7zmPNa5lO2uvU3SeqCa9oIosfXi/VSkeV4WkXgIt5hIzwfPd1bL/4PmgcTRyWuInBZv
1rIEUdN5oN41YghVj+xyh8Lj1D8vktCWpV4PXfv/BsNUZOdr/uILrjYuslvql2/5yS7vDa5eTHlR
YG7DH6IkoEMa3Cd7cTnpJ9UvZilE2xEn3IBGFaKd2WJLGnlngLIk9Brq+XRc38WPzu69Fr/Lm53+
C6SVwxvr/Fe+NuvzMiEewoVw29iMBzDPLidyysrNog5WmzXHVqe2hcSqo7Js6GhmlSFRlUXppjgY
/9srEe1l5Yyj9UFvNIca+ury0uOaO0K7/kz7D5+1YSLVQh/JZzVMeeKwt/oMEtCNBOVcLZ5Gc3y/
kDrpfvgp4BwKAvhRVSvyfla1UofqWCbfMZm7h1wHoMp5f6P28hbWXbnZBCXW6yIG1A0ElgZqa6ef
LCDa5Y7VHFgymyMPetXn9191daYOuEbsN148L8+v/TIY8dRxI0GVjVTFe74PNrtPgSAhYdTtAAYZ
708yMyNTL9ckKVIDc83WJunYUj72S1ARWdCY06t6MxOB/TtsG7i6wSEuct9Wz+yTlHBDRyfznUM9
tQkBEGDvGV+fo/+JDuiZNMdY3Ack12XGY1IPYhcUuyp0sirYiEtyum1T58984KVUxdv81kxFRIcD
D+g20qIVbCQ5ycrAd1IdYHhLS/PvhPhPnP3gVa8FTSK8KmLRWNdedPL7EPuOdD3xOv0e+wDl4la9
PFpb02UjoaQaCY+oR3LyY/Izd3OmjkjSFpWMs1eEkFvhvJ7DmbixbkiMSko10PgwNNQ7m76wqMK/
vWGzho+1GPIiguCMK27LwlUWaqV0UAK9GB5yEmbQCLuJkIAfGoXTJ6nZnqz0i3lCykIOtSC+w2dx
6h+uq9foQc4cJbp8PtJRHCPWZluan9N8jWCsMYAdO1Smp8gJOB6RdqMLC6bj80o3BI9dbH2/wnmb
bpHsATq1wpFrRQNUE1DkYshqMsltkl2vZ8mhE/555yKXuOpIa7evX5gQWTDEQqNTTFxOpZCQZ64x
iNOEhj4RJ9eVWgZciR5UTVZC1puXRas2KAKTfmh/OVtufWOGCFmsez+/KoQS+XmJy0uPe2J9TA8w
SPFipAn4zW/QPIhKKaY9cmf3hmbne+mcQx9DE2/j2mEorTP8QufGH2b/+DeAG4cKW+nJau1ujytJ
ppraDAyNC3sZxLaqTOll0XT9vsyyCRLZp7F9DAWyj+FRTE9ZBbClQTgorN6Oj3ep4v1zvQncfsRZ
EJDMqaUvd13gPQkgCrceg/BQFv97wQs1pne8Rpm6vy3hrPJrobxhB1atx5QhRfbE2+7TIo/BJQe4
TTiioaHvH4QeAzxI8wPb/6Nlj/vJfVBAoJLmrNw1tgNcBN/BHDO7B3Y9W1xR2MZOOf5e3cz4gwT4
A4n/YqFnWUuiuHTmUKphitOH2CAWxB20IYpY2HZkW3jLIfv/zZi1RHN2rSTUtqDme77GzcgpHhkE
vbBW64BRNhN7Wlu+r5JetzwVNxRIEJ0POy3UslRIPsclbeKH7EZCSY3NLZFbPqEk3wHryzaDN0jE
fwCJORsGsve71kRNbqb5ESbhEMFWgsubOxTSb66UL9mXcayt6Dg0ba+B5sngquG29H3TyyPtca14
Q9GicAXhXaHn8kt4UnY+VhefYLOm6kx6+Qn7lXse/HpMjRIG/1p95eZ8aaBwctY16BiumcOrNiKA
6hx0ZD0dglxAASwN9UjjO9RMxI8JSyWt6Vu9+h7ZFSD30UrFN2WKXiEHBMmx6+BdHVXBkghajFMz
DJX6DRLy9lQTSQbUPUJ/YTqUf2NHp4JdI8imr0KEpX9kunEd/y2NhcazXV8DjJ1xXNOIZGOcHbOq
etWl3EpEQgfWn+326msE568AwSw3GKK2jkqAprOxsCYry/dEjKgUsBIdfLua1hBtJ8Pt29vQD1Y4
rCmoqsr6VQn3Aal25DNOkSInMdtf2qppx7H04+/68dsdJUQ0+fPpER902jVKS1RuV/sP8XNbSQDh
3oW6RNdfiC+zY90Oso0Gm+Q2sGcAscW30ihLKuDWn+wknRuUDu3wd1idKX3MRaqmkSVWrlkXy2im
go5UlVmHMUSVZF88isl11Q6t55XfGIA8oZ3cDPtxo2op+yhlAXU2U80OCYhTPkKrw4RnA2mc51gR
g35rn4PyBdVqT6sz4X9F1aRHfd58hCGbK3SYlmlE6Np6PtGBzLRX03NNsHqD+VaUvJ183Bz0hvlj
c6IkTMuwT8leZLsbMVgx9pH+C2nmS8rWEjgmGbFb3TITyemhmZ4kqdmLBXPt1A/Wvhg31zOLDoN2
L13YMRUYwJMjzdvbdWTOZ0nSvPvB4xGHnICAxm+cTmhFADaUHr4R0dEvs4c95qjxxWRs3L/8n6Zg
CS6+PqmfCU5Fe6TB6Y2TMPZdfORSNssHHzMy1r9nLG5Og7GaZUqi2pL7DvJtymPAD8Kh6+3Mu6LC
Aqr16EKVlTDzNMLA0J3AYfAUYncL6yXFMThoSZCYRKGLK+hQCUnx28oDXKvovcs07yMv89Qg1THp
5jz6cNYnq1PsyX2X2hdXmlB245en/wLTKlaVhK9byIz8UGWnQGc0Y2slXYn1KrdaCaEQrPRF4fz+
nPPvSMxMhn+5Wo7W5KaMLuDNgARFHNLG2i9oB1eru6VCi8HHr7WWkkoh0iVtAtjAcImNJc5b0+f3
WeLyAiRmcZ1wb2idWag1DjHCQNJEE1srpyJXft/lg9nxCO47b5ljmNFw3yMWnVgsfbWdjPe+OeTy
GY82IE8ciCKQi9MKTBYhg0T+En8Pbs5i8bpLsImLIH+bcLG+13oF5EgPmKQljuzIPi6RqlcCMaLn
ZDKSgPLfCBr43ZSW8tWZvkvnZmfQgouIRX4SmMf7x5vfoOP1fyPQukuiqNofaw8MqDQosJH8I5qB
Q2vTr45/Ub8YC1IkLRXlg0sXyc2QRnXqeQpyjze4enrSDLAwggS1QIfbVOa7eoM+Q9gXyMUrZoky
omOlVfeWX45P3gWW1KqBBDfV2ogumitu79e4B9KoLG2wFmOPmMte54qYUojWY1flJ5uTCxfnFfEl
u7hFvBBUxvn8FxqU9/lD3QIdCfoJr55BOeAGQxZSCqEF4xGCFRGBuMBVxkaOyMNvC/3GxbUxwYDE
gtxqSU3rrMtelGkTgUfGFFEmiiiT8jAEDJsQ3iOz5h1MckdxY6+DhTT5orFll12D1xniiVyZPTrF
RlAqGLIEcELFGVOTMyA/vbXGPwLB1iC9VPVPs4yr1e49W6+lsVIhPIfQ52+c6QgBCFJsbQ+Sz8yc
xlYQTrKQMVGBBhWoZmKG95ySv9ljBqSjelJ719eZm0F358e+emCewCjlEDuoeJdUeWVCTU+eSf8T
wcooWIXSrDbBTdb4DETwaadSiD6zGTo0tH3S+ofiAKlCkRLs7zqMFDPScc5QK6O15LLSGbwXrcNb
qNqA7Vgw1J03vHNtXBNN1xh6oJ/U9Vb+ngxyseoOqr4NGcX892PMrMOXvSj/cTsLWagyAWY6tk1G
y2KBpEPMCLOifBN0PfuxPaPand9TOS+gBk0+mHY+VmGOm89H6uhugmDb1+NwcGAHeIlx9JBnpAxq
3WfalxCjpy3EsstmNKvwT+0Amw50CsT506EvnQT7igc4amrBNIvgpc0qD+Avz/bkNNswxzNe1hot
MlBzXUBolGEPZg1wrtK62wczbIHFJIT/WSmBr8prdSf82AD9BBfQlm6JI/QdvMPN4jZ0vwWyi9pW
YVwDAryWctS9ptJJnrTk3iPx1Vul6AxvqoJU13u3WlNAroDcmWezcNEmffG8MVi5/QYU1Ie/GM1/
aaUBkpsCIBo3waVfO9z0QGBZbefP4kp6wR6oSrZJic4lPGbmjClnQN2Z+9Q8oSzlAb6bYYm47DTW
/VAUsRFguGDC5IDATi+CXT4sZLz0JvqsHODACfLcgTOaNF6coqfU3kwXLJX0x8EZcQHl7Pzqha9u
yiQyhmPAxgTFaA8WaPjsZQGcWaW+wKAWVVQilTbEu+T2kFQsZOVYIa8GcgiGkferhwfn45lLk9PH
LccC3C+hN4HByBiWhGzQXer9aIaJUeaOLTdOBBvJg74sPvrtVd5zRiZOgHibXtHllmNRIMYnPj0y
HyxUHun4vytx/yyj4WDn3sHFxmG71til1eZilMxuHhCjiAZYuq70pm/JlR6VvHm5aUODOGNxBrHl
4aGBLANprKsfc39w2/Yw4I8fnt49Tix/bYRJieM8t2GXoKcPwjGNA7kkF/cs6JIu0Z6Qr1ijn2J1
f9iuy3ntNHmQEQildqZUEFPYpBL4dL6CDgiGRNOCkCF4wVPZTV0B2wvbKKSL79C4lVOUq+qhZ2ZH
ojO27ZJA6YUWGaiCYINajc7r33we+X3Gz3GwES8xv+8MfElV1ZYxZ2XSo27R4M0mFHqhxsYMw9Ir
iwWw5POGutc7hJf2RO+ic7MBLkLJwRX8iZQEmtj3gBNnLNxHF54/ClHR6DIZOhRtw8drjNgAXeuq
gWQf66LZbqN4uETFUgGqyR4t9Omm4V9lS1JpwYaLmwVcUK3vV9AJcwRKowCxWOf5jLBz/R9IV1w3
GJ3fHPNMSIlaget9d5xaQWLVnzIYCLAfDkg34Osi5x8Izu/MoQgOr1D0fTXjSIcz6vyCDfGOMXSa
vvJNMUjISOurhjrd13d6DFA1SIXh0dW0uP5Nfmm5L45gzJ1ZyBoKUC2niggHHF6CQ/Z9mwwDbsvP
XbsRVzC/Ilj1Isx31GRfBibIGZAoGamRYvZL/LCjd+kIiIKmJKAD5irNTHTt4Zb7ayXqO9J3bGFP
KqVRS4qgHED9Oyav93qTomOLZX0Cz8TwAMVAft16kEiUAJDQSA/QV8dHTGC9y3LD5GguUD/ByNhi
DGbAUy9hronqI954NJ14e5rAlmfL6y0X8Hsem6RW1xHu2ljrkl4YHelfTzLXRrCaAkK+wVhcElOn
q7iKvusAtdFJeIYR5O0ptXjrkFB/K3eLdmMm9qiy7apyqECx5NObROUt7NYKMAsSIGFjiIPsgx4M
5EUQ2Vxr3bUkcvpKLjgj1nSzw+eySz6rQrolTU9X+xiLUYCxQUDu1UfErMpPqcBuVc57wEbhTx0o
dlhnl+AtxLRcjvjwmkE5ldM3YvJEtWnkqgeKOt8+DF2LqZOBYeuBw1PcqIm/RFqL1vgCqhjY65v9
WuQZ302seTXULIXpQdcdnoeYr8J0SigAu9RqVaBeZJ1j4i6Loh/XdVTslS9PGFLcR8YDBV8QKycS
dn55F6ene2m4ut8tX0BZT15sXABP5M1RXTqxCxZW1RpaxQdHhMn2QkpPSZuORQOUlffedqa2ownu
j69IiLXqXkRoMk6Jzh6+lVmw6HyxwgvLgmUHH5yIEEocM5T2wo33utvDQSS6mfRXQRCRxY6zHKNF
EPk2l9SD5kvRXaj0dJfC+sbwtcBUXYdj/DEF0zgzxafWfyIbW8MTlXepL0mzQCQOvNgQ5W8CgbAP
xJyNbtQR6/UzaKBdqZaxAHkmcGgm+sV8yhNYX6++9g7wHUk8LRdPkvvkmCEFHkuXPijoKY3mGh6c
8lnMFq2BeI/PBfsHe+o66GLroNwzRxhq5Fj0FaL5CTledDttNBfFT9AYYB6gEnwdfyw6zcVwfyci
cra/4f5TJWr6ldNd9UxJOW/ISqndhCl6rRWEyFrTrkVVh5P4ZU6KeVlXAmzPFWOsxzlajJ7TjhhO
nHuuP600L4zHqBsL184o7Jt3bQNQS61bWP7zuLdCmGtaq2FXSbz3PhNqkUA2haeuIIXhstVbDLOR
HLWkZJYul3SG3a4l0y8TaCdfUn1Y1sq/fjzOyN5oMZpA70HsVQPtt8DM6D3wsC7T/1WsgAknhuXx
0y+41/ad+vxixf2yk3D7iBylfXZzJJp/VZgtOvalISL7QQfp5X6VSAIHMNrY9mK1NUvOQvDEczyU
6kpNLwAR+j6Xm6dSNbX8IxeCrPzMoueW3U9B760zGjsAMho21pI+ur050XLvrruSgA0wG3WCDMro
3myE3uEm+eHJI2AppxtBvss97LFiC4JPv+Y4TyMD9qm10ixHthcvWekU1b8ov7nT9Htln7muMBT7
M0q+H6bnvd+XvXQqdSWJ9QnlCc0YWL1hPtGQcIPEcCtD8W+ywKLTWviJEFVvcgoBn3X8x6euUENy
Nbe2sdyNGFsM/kcQsUqlm3Qu5XK8YZ092ey+c2VFUalckKkJsHw56ADG7qGaA/Dv2b4BQpto7fdW
yhWwNdxEr5OOiOus1iB/ALu71Gh29PqcRehYAPetWDMm3Lret3dfDz64pg+7f8MDeZATHpsqkExl
7XSU9Ytq+lN1jIemkRlao40mzQydhh9zK/g2zxRfBfAUcDa9+JJNpCKxBguAROMRV2FU+00HdBCB
6kbnFEXLKdiJckuaRMmIudofvbv2McKPZpU0L2VJkM0x7ThHs39ihRNUbwUNt3U2fKdqfAwCCDxP
WvQVwsRfMGwaYg1wH8wc738C3Zbi274PffN04efU0aH334ICszkiJla6Nz4byxt6l5oBztorPncx
SeuuxASIYwZMNkTc7I1ENDLGCYDhcTzxnwFTObP23igYAB+JYYzFFfXQWdo3u94ZYRY4FZs2Zv68
zq87P7CQtgn8m9nNv1KzfSI6Uq0tFpTFlvNS1Rmgr81KMtutuZKWMcSsat7jH3uq6mBVOmUFC/Jk
RqtK7iGXmTro0Sf02FmDRI0jj6unbuIiAnooRIHIm/OV5Zx7fz6QkgCj5/EQyKlKfB6PxMmm/kmo
0ps+7HnfyBHBq3EEhRzHMJscaMNNXIcCPTdpJmB/PDq9HhKEx+a9V9Q/0vboaXYd66tvziWP+XV3
pgaqKKtpZ3/t9j7WsqnC5Rst/GnMqtFfg9m8kmGiVU/8B+s2UciVTEShnCaFD0Ro/T3IBqGzNhAG
Q9N7lUsq0n2hQdqdZrCtqf3ULVBYZUefIyDHXjsrZfdbdBeMtnEegem8dJVvhrNyU8L/DWIKL5v+
rVwY7i8BYneykz7YtuP3iMVjEjzuBumzfH2Vk3mZfBlSVx4a+KxwDY+BjbAtNHiFtyGGlhB0C44k
3DnpMU4VWTh1deVrCU121MwNTFwn8NIVN8vZa8jfVjEmkPKl7eImYw/MTUsdTyXbX6nxPxiQl53Z
XM8g/k8Oy8v2Vgw3+z5ZUg476FN6cX2exy9Ejt77wdUfJ+nXVibhdWz5hhZwwqTEI3t/oKAukAaq
3zFWLIVZyf/KMKdFCDtUZDZNZpcnHFA4r2ovk8WeLcPaAWJb6FOElUXZN82jBVyAecdkSTKB4Fzx
ug1L8HA7NFIzdJ3lPOmE4IxYeXDPn39DrskLo9L3+jMZI+Sdk/Wwyg1E39/5AWWN8/zgnzzeisR7
T2AgxnwUo4VXKSvV3vwaNvsFzLHpF3ECrxcMbGWZNCs17voAApM0oY1cpc8HEsEbjw/DlyH8SNJj
fPPs+nNEhcmaUadLEnsSVmVehvA2VZ2ci7BC6HVLjwlCJ9kDjC+fAnj+oEEBon4oj9qZogaxnojy
aABtibDTd8ma0HGvqHrZbxAS6lMdlxyLE29HqG8a7ZU9zgfRRGQbIKG4i3I/w+ItpRqV8PxUJFzl
g2lS+NZ1TZRyOKMEN++PPwgUGmo/m3n4RPUDRWZoev0ngJWWH7E2k8a2YfODjeEcGc5KoOVR6/FD
abPjlVCbO7BIhB1IhL/Q5OEHZ88XfGC11l7GUUGUxi1TjBOzpWf1CLNfGpyJBBPULCK+bsNxVfVK
4tsaPSXrgeW+BTHDSD9e+0p0LHdSXjqHONHBgeHss30gHic0bkIYTW1Iu7yAYwORX4kvQMfE569D
cCRH79l6D35MF4h3dDX9c0wa2r6dtzdoumzD2tCkIWb99QXZlxaooU/xVvDc+ds5S1ZSXpF57f4F
bHv9pouX40uVQz2t6zFheAwM0uZChOHqO4l8uA+10GNl/LOdaG8kG2RpzL1DU7KO7ssjegWzvh7s
OvwCQmV8eaw5nFrPXBya2Qx2liHDf0NXlZgsDjsUxF4r1H/FXr8oyuU4X77gNHZ+2LLcNh40rKjj
ON7W6EU0OWEoiJz9mypzyQmklq0CqfWp0QBEzhMQPhFCX53QaTiUnuU/C6zTP4WS9XAg9nF8H6RB
Zix6Ttjlgp6VOEpFb7AuHimC6bN8eGUqGlBqC2oHEywYorU5ayOdcS2Xz/me4U0ir+UauiYrAPSx
eRc9vgedqOCSFR0p+15Ws7O2/ZXfUxHLC1zFnAXyeBa1+6lA0oO3bbBzjwS8EH1Yf3+AsPyBreFO
4O2LDwCj4lRl1G6wn6jbg2nD1+tDHPiUos1TeJLhnq/g8v6GX1egpPxrvpGNl8J/mP5KTNF0GZo2
wjjEJnWpueSCT/N9V8fjwC2CqU+2qLMRQU1l8rdty/Gdl8HXx5sE5NlazZkecVa5DuvOHP+AZYhZ
gKb39nRgtE5ynGOKxaRvh4Ees5/97nlkWxabgq+Wk2DyXzzEvfDL7BEArWswX5nDz2HRCKY1tUmK
/3pb04MJdY9TsGvltPBaoByfh+r6J1y1NOFesXS0J7C2Cxp490K7m7B5LhiSt82EN9g0RtPe2CvQ
ATKwWRXOuT/r1YMXza5VjaoyL+Lr8q8I7ngZAVcv4Znezv9Eav6jYvqjQgy4LTA/5dsmAd6ZYWVD
9J+L0QEvzNWxTno2E9E0nzH8ZUx4WVyl+8xgqwqHTSu9PxBj5JiXoxUuPkBOZfd9JTT8DDF8yLZi
1yLTfw/xhEvK0kcqMAtPhkY+uE8SAaYPxGTn1B+UnUQz0+YKbkbiFolILMOW5chM+BsiSALNIqBy
cu7YRVsATtgQ+NidK63xTOxqfRzY49KArQQh0HITeLR+2d4Xmm84TfabYGfQsLzJRG5KGLNZa2vT
NC03ubFt1AXNEj2YVMeDSu9oVmEy7/aCnw1Fpe5tCKdaOIIKOMJNxtn28yAhf+zYdXBo/uGYjGz5
kkr/a957EQM3wkCusjxS2vxKo8todhdkMDXOXZWAgKmthR5oquiwmP6f4eEtvb50vjkIaOxtN8SO
DxAM7MzVSSGQTmQQsOzoWGynNVDmZ9gXP2xHTZdDOCwZ3fiq0B+oOHlbkffmEICtNdUE5F+EvM85
fSW9sY4/TVqtXtkUZ8XQ7gIAyYLqwXqNn9iad2M3ipiSzl6Y9z0/XmMoRhf4XSDXaAHBe5pcA6MI
zScvNRit4i/qvS3Ts9aqo69j6BLzBo+6GAfjyO+kI8EDXNT+RRnRDwUJ5066ImOeoMQgDDZBmC1l
ZXiYlzcdP0rqbgZND9VK+1+GIiieUasQah9fh8n06d56XAg5Wcp4FdBm4S2WsumwHJN1w6CvPWH0
x4HL1UEx7D3J/yQ954GtOEa8KYxzpjBBDzUn3mFa6uUV4kEA6R59qg/XVDWjpJqDcxoDTD7LJFdt
RliislLqskiNQBwqVFLw7Y78jeGssgXJOd1uv68X/SA8gt4EuRILLSFa76HbQTydxT425N0c1x71
9Yck4FRKV8FfhnBmmPbl8PpSgOjYgnAxXwccdg3xM5zVcegRMG0Q0jNgyCQcoil+O4KC4399sjJF
xvghr+RchvUpovstRxMdnuoiU+GKfYN+ftzrUIA0yxQYGWDvHffNTrGK4sH6vpEb6/99wNu3ht7g
Vz16F6eISORQsBQdoR9BvNXBnkDhAInZSrTvTUt0DLIDDw/lM8aG5pSaRVhsMnyMHkM7uVsim8cx
Sa1GeosFaY6+Lg56r/Xl1Ch7vJlQMXFKN5TV76w7uMlvxVFXV8oVJe1dAA3VuPJBzhx+5dPGOtdr
BpAbbGJkH0t8qRC8juNe2Rp9Dqf2TZhaK8CVWpn2q3oX9MOPRqm1JZeV0/e2P9eOu1ofLKfQT4Cw
0xmWC3aS/cYzNdvkVuRLlkJhy2zcIfXTQ0qphOucxGKvf0rU0HG3kAlBCTvCyUnb2CcWmO0HK4G2
AP/FlV6sPKhYcznq41Ok8ifIwhqa+Uv5JQSDa7Yb1/bLcegkU5dDDDVotRqNDw4oAwB90uYlZai7
DVzf+yTSaGOJZzTcIg146Hb6GBMzGi/zwHwmMv1JCBfIPNQrGOg4PzJehTnwn03l4SVh7YEOyNJV
Afnob60I0mo0ZZFckx5ijswW1BbKut3O4bvuIFCFrTiuXkBSYYKZ3YF5Od6Sb4xQVUVCIGfZaNW9
PEU6NJP119+S7yvvHBsBplNF5Em/6yjhUELsv16CHz2juHk3ECxvRkQ36JJ9PRIEylbt7NPJl5yy
FAuDw8vw/0xd2kfs2h0yVIGceGNIPVfuazyqeCVH7aoj0hI2Qo8e8pqPT+5zNzhUBDQP2135SO1u
vDoTuos8x9V6nYyTjWHdkKVID49UTJESIeZ1WoagUsV+y4WU/r+1LlmjrwP/yM54LRCfW1FrL56f
5TIwzBskvKRUga2U16zTGqPMtSqA28C4TMNdJhuNsjz6BjP/9B+HmtU1fsKTDE9c/jQQdhcQ8Qcm
d3GQJLxmiYByRQaZNn5o6XlPHdVGhFPdi5IVh1LcScD9bpqwegYZYmS8J/B72M7/rNm4+l6S61lO
TetQQc1nWKpwKroq8h+FLuTvXGtIZsbHFDwJYMnzta3UhTrXdBN5V4egX/sOIpvWe16w/6lcQE2p
XHWBuPN/LXeEN1CV1xximWJxFzICWEGgqlUI9GdqwpD7lF9RQj49qmpK04w6UX1W5Mkipia8TDBH
5hyLoJ1itlJ10KAUmF2O3Fku3FXm4xw+pR6npElZDGNdI7Ww8/9X1SNMrto/uzRbYUy9OjRASXsA
i0aoKa8k4krS7ZnSj/QJwZC+XchgH/UyX7L3iDCNFiMXprgaForZWHXH+k88faqCdaXUHjYVLzcw
l65oKC4JYx515O652CPtCmFcjUVvI0uFvPZV+/uhYEMbWrp2DG4CYmt0A0GzlCUFm8G2Gh1TOoCV
3K4miKa4GCggqMGJSjrPUGvC6Q2d17MDFzqIjR9CThNTIDm/kHXTtWAtadvknKxZahCH0x47Yevs
DoJGP/IZihSox+sGo8a03cCUn0FJsKUbVKSdyolZwEsz2yBxQQGZgNJ8OffyoRc+IdSU8tPWQ9qS
PskL4hoVssk47rTraOU3itrn8/CMFUBhv0aLCVRTg+Hl4+fiiyJVP0eLpjzyqn4SOGQuAlnu8hgS
LQcJdcD2wkHQ4tiNgnYJryYjVGc0n0BdqJfvtE26Sa6rrrW6DpwVZhfeXK3i7T6sd1TvR3CK1LQ+
rnevqhCbD8D0YgCe+nJBg6bR7tR60KEc7IKqFHYzBx7vgb/Wqu/fQ+KG87dMSoXxE/FNnTS4BZJv
U0EYNboQmxZW9qo8JxNZO07v/UcZzfZYbRvSGSjxKBohrPyqlejIPPx+h/5A3bK6pK3yQb3J/G8L
1kbsPqFD8pGyGqutxU8q5VvxCwekIvecnjI8Zn+q4oNNvsNJM9wfdreYDVfBc7vYyd6+JMeYXxyT
LnxRSD5FT6J13G/Uyqbh50XrCfR/i1f6ma0j0iGjIU4CBF9gmNHV3FReKYiouiZbWF73Go0jXiMj
ZzsYOmchw+47Hwcen5aEZZnUmR0r/yqAZt+S+UplI451Ah6UdNAz3avxKNEkHPU4jlwxJKyw88od
tFybvNyw8e68OfXgp4SZoAeLc/whr95nsVWg+YYGhoXRtEZPWUghntfA635AGL+crROViFtzlZyK
grcvlZw//hEa2SixQ2DhvFfHoY80g4ypemawDR1GN5RJxN2yKd0QtJcpw3nUEoxyZhsoIJ1uKD+A
iWCb9LqmwILcIAza1BpszK8PIqMtsUyv/Cwv+U31au0eaBcHY6xLtBKG2+QoXXOeq7V5M6z8jD0U
8txYL/8za+b5dvURYVtEA7keHJD7/CtDX68OeIdFQxVyYAlezEIbjiVW9EBkJNbMgaJngUf6yhn3
MrAI6TKpYCEaVKuI7uPbPb83YfUm6mP7vRC+Su3qvJSlargJcrF0QGfsyw1SHV1t/gtgPNjfU/if
zobk4XnGkh/XwHoFo/aEVhl/p/OGYr6xA7Slr9ppCEXkw44ioWCjqLRrw5hMVVOP5mikyEMNsVtJ
jYAQn7w/zL8DpGFN0MUBseCaZQJP6yvTiuer6veXlzIoyaaTmZZd+vusw1/qy5ZQJCW4MJaLdVVn
cTminissXRn1fm3GzsCGG7VN1QQ/ZcqwGwdpYrnIJr2pgJUn3/nMIsW2/A42BrQSxd40xcnuuF+W
Xxa2/89KfmWiCt+rLrlyvQ4emDVL02AqxO3cY/BzN7RHNx4pC/j4AMa4D/8rBBP1lz2wlWlQgKaG
4LUDa+XGNeD2dACNzqK2mmNbFDfAM2uq36g7tcUErJN65b6wiCwHDKAKsKsrhfezspRX1HLTRYFA
4RAbTxMQG9FND4g0/eERkfqXLN2LfWj50L8DEJpLD/rKIqNPG4oJwr4dc+7cAw0R9gjxDYoPbPU/
bdTautZn6oKh/L08MiQNBjqYE3xGm9r3l5K8xDLDBWebXSIQ13d0mreg1Z9laczek3eq8eG4vcJc
K37pr9DAsju1KLV60zVDuDievcJrOBxig6gCiAFvlDKQNpiJ/nbI70pnNOxUyVVzN1K9RM2DBxh5
EysfemwKk/QC/09C5WTCS/aYuXNjyhHE72c701DoTSsqbE4KYTgAtXOePTPmgAoJjDM82v3GTeyY
3zD603FS5QfZ06Og+nqg+wKDUA1AgqZWzIPmpVCT3IY9M6NaZ9yddFHwfKvAoTjAAHUBGcPJChfs
0QaYmXgZByAUo6feH8xMI+75A2kJBGwq3b8PEmxyHAfKh4ZsGYkCEejcVny3POVJrnPZ2SMGloxU
RFwMFd/LeIU6re43/ioR/WRBYgyYq3u8hKz3mqoGzs3txHkiSejEzb1JlXGXyJVIcX7edejI37wF
mRbCSak3f4fLUOKs1bNyTmZ6VKNBI0yssW3mDiWPX629QQeFcLVcS9S7Ck/DaghcUR9MY1j9lFqK
JxS5hOkWvgm9JQkkUKgpEq/phl4hPIJtEtU6oScNeolDWU2xVeX1IbcRo031vEhDDkPHwpzPb1G7
yr5DkK8rRL7Q/InqCIpiymSJh1DlAi5s0GhNIjxZgDrtKoOhVZuKWAOiCBtr3KscEUqHSVMmOf3A
W47QRIqFyGlhgkYt6TkpMK42LNsMcI7tRmn6hr7a+WF3jH39fY3DOvd+r6cUe76F752OQWsFk69+
mJxE2JBo2YOu1vDkUCI0ZTuSzP9C/Sgipkr4sU8rhG76FCjl4ExD3UI1cErK+LarDEe+qrvQ5Z0h
FQQ8uUC1jxn3n/Tgfbx77FhqEbs8JBlrS8jrB1SoZqxRJuu986m5ED9LFoxtqhg1GPH6OWrIRS5a
sKWBGWp7Xxo8sHd13Mgj4ozj7h6RLYGR88klIqra49d8G0jTJS5q1OUQjMJ2XQ+3O0if5WJih6BP
uEKhHmT0U4z80fXH8/yKSpQilhDB/pESIceeYE/e7sYrK97gw0ZadPUWxGnvfJOG4Crs6SFMHvUU
skJx/4Cf+X6Yzpg1su+AO6YKU1pOnNp6Qti8zLRA+Jyell9YOmJwpuJVIPkHRXEcfhvAf0e9H7V1
B7mUXECXGbAQSoZCgD69rHZ0wiHU4tunbaRHN3cP6b1mVMtYN4MB3CFoWonM+0akCwmRTc9FSDXb
OaiVrU9FzoIIWWmWCFXa+aX+H5M1K0UzBIAqgaluQqpxgtAP7HH9h8ju25bhRGLAzWtdiMT0RDu7
H3ARO/Z5DG/9aergEKkFMVJ88dYC4t1dAI/2fut0s5EPINQ80+ycoYGMeH3zHLnJnxSJcA/VDmGd
VV2BGv3DwZP+Wwn7i5Fdl5uM9AghdmuAqZwLKJs5v0Dh4/TBOTVf+3EJUVu/uv5Jyy1uShVX+HpO
UiGE85G7GLQJTmnFBIKID8EaJj6nhwYvJpykgfijShal6bmgxUSEaekEOBl+os6aCEKE02CFtFK9
1xWeafZWkS1FPZdAuutuqydDXKpGrPwpXOQWs1uKn9745YczkC7Ktmr6WzHjKYwSaevs/TNjwnfP
4vNRg4v8i9IbOQq6aD0zJoRT73KKUwPagAFHljTyHfWk3E9xH0Q77N3QGxkD6zy2lyQPCOfkjZf0
Y09Oga6C1RkKOWJ6vTmEjH+DXy1eUMds8ogEF8siWfcQjPnd+1JXi2ShCGkK1yzDhTj00RBYQvsM
KXLtZtkH5KIAjcamDrGB1Ui/UqeGuDiD8cUieQ0UOO2nWTNDiq+CjELXFOHE9mFt324DPGYN3I8P
NOCT5EOitsny5+4hNJU5A1OgKHC9+uN+PP+Al3AEyJKjgIusHIeSMsEtFeI9P4IqRbk/omxoOy5i
X4kmnesQJF3IDl4OWNKqPWP4/Fs7qPTQXGBMB31MaM3dN+QZPcLYZhs9ldtNMVYycwsza+00SvVc
F/Kwryqeis+hFipp1Updlz7XB3hqaNlSJ6PrSSEVY1d6ajNbgSBjseP1LffEGJNgMI8vyCVQlruX
sDqrBDOwR6a7KFTtMhQTN/TRw+GFmWTy2bJB/KTH6U1F9xuG1fHwLDxWTEU5iyjgbedWcREfq12n
bRNW1O8imzZ+3WdU7g1xZTjsRzuu5+nVWldAUMbnUto9kjoXOoBu9Zkr/a7QOupYFC4PSJGGLzEo
hXf0RMVF0jyehGfxb3QyH66GKhT3GKQ9qPFSrSQoeWWljgZwPXaSuy/lfMZxKBcLtoYhdYm2rt6g
Pkr0WcwyeMad4fsm6YJ7ZvMmLmkmaNPBoIQuSMqLOoxmX8wIqpmoq1k0q54AYvCwTElKsTvYW4nh
xbM4hAEAenKojS/AUbt335tEPALBnC16FkkuvBDP502CIr5DYA1JGJkuU7C9HRrlMKvy8z5Ap8bv
rnv3g3JbqNojGHQpwZxdcpAcWKI7TAcUEyJHoA5H9D/fs583KTy4it0gw4nGT8oGqAdWwN6r4/vE
pBqtb6JcQMYX0EnTYxdhIdqhTZfN91+MgDh8N33rADQBI3TfvY7P6ZQDg8vMIxdyZKdc0ClxcJwi
gzH9Gec3lMWpMbDnNv9LKz42JH0aNl1DydNETVQsCnl7JG1PhhRb/jr4rgUxM5f2QHpB8b3bEtjS
T7XzByXYiM6UtKORGyC6iAImoQM9yt7VC0C/WVQ/Wx/wkriydVp8WkWGda5BPh2rT1iku5H7ogvy
/EJAYkrY+OwrENRTCwqA6cGNizjJaeByU+y/cU8BJIfquqngdZA4NbUVJNskRFpL+Frq2hCQjB4c
vLEop/oAdw/sjz5UaJUJRZtl3D6d5DB3S+y6ybNwwt820ChIexriWM3fjXMNvVQyZMkIEeIGnpjp
GiiW5dncp7GShZgLrZigK8IeYmGEKfnq5vvPjS5K+hVrvH3kKpmWsLXaWuI/CETCV5D0gKlBOyoX
2QuuV8ijkUmXZt7YcCEFcYiHsDu43K8QyGF8xj8ZgUBPTRFJJU5uWOda7VabRLXefaWF768dzTIl
QiFGc/dmBFiMNdSjdLcmD/1PzuuyYczE6mQqjoRckEDvB1/9f7fbrmPB3kiAoOrBdgmRez5JkeqF
QumyZFVAMLHtehh574Q81MQCUq4mTsqljwk7DvUmeFvXNCgWBHUJQ5T3wjCLyyeBdudHVkblYcz/
jtvvfA00O6/zPfJx52DGI3LeyOJlbH6evJsg1HBzloSdjuPp3SlRWMWSh6naf/+M3z/ASLEzo0cu
VK9ba0h4mAEJGdUVdAXvG6GurhYDN6YkZZUA5De8NGiQcTGcsemzBu/KrEznqFpOExmNhi2mgHAr
gI8n8Bdw7z+hg2woOKx8hDsHHTVfM85nxhnbuDBEzVJ5K28/FcyqS2Nwsv+uNldnliasw1YQDDax
A2dd4Zww2mhx6uhM4be7vdu61GBNx0V0Z8Qp4mmayKVOkEpdnWL2sJfAldFaAcKQzjAQqRIAmqEo
5E7lmIom6885dBEdpo39jnbcS3/x5dZjgkEu86TbSTIJeX1VrwD4ks/nScZ+lMlwjY+Lhh1MgaQ2
1K6lOzjvlLKy6PO5zLR1X8ixzl/+cRVRchfFZ5IR2PU5yN2auqIaEKJLMCyHVoIErR7O3Qt9kk8a
SkgGlquln/hhUkqgcR0xT9aWBRy/+lIvzhXFVOf4WeDqAQLKg7Bw4Eim7X/lVP+LiJxQkbqFTeQy
QYyvHOyrs58TO6Id2pNsq/gVbFi081LhoppEYi5MaqA9bl6+QDMAg+BQGMKeCExY26+2ASqjrbIa
ycCikWlaHgWTGu8jkBQ0qRsBoxc7V5GEjNKNHoeL2fgQIjatX3Wfof7O5wcfv6LIO7c+z8DsfV60
HcpYlNbJ+RfIC1o+XXiSwuTtnAyriuFIq/qna9e3nEc2dJ2RotmearrV/S1S9BMxoYUVBVb6jWF6
/QvtUx+Jak7OYnbVtpFk0VWbUEWfvBn7MF1TGRwdxwmtxEUgXT7P3vbLZnxh7helqEtE6qBqqrZK
3Hi+cEWo9jgOsEgphVgRd1HbQ0DTlRd7F6jtp/OJeoK0Zy7uZA5d7klivz6x4OpnGB06gLQHEIww
awSNY2ODu6+X3JSB7YBOURfrLakz/hLaItIzWC0M2SS0QWeWGUo73CdwV21PFhRiKEVG6RUYxWuY
CE1QxaEEifDbM5sodH7Ttv2TLpQbw7O+mBE5icYfAP97dwBVVPk1NZ1TgJHYKERPXlsyfzQ1rFeg
xO4IADRnjf9ewfFWJod8h9wu8I7qitGnqXzHxjodM66Z6tLGLMOJZPY4RI1EUzQ7fLMGPBf3BJx2
UVXgYY8uvq8UoaA5BggTwqCupCOSwt4vz7QP/1DnwQ/bIFDidkJJN+WXVBFgjQMrPDoye2DnNfZT
KjqGqw5MaPvebnkfp2R6AOcEQfHDxhXHneDua2TjGyMbqqVtxpA4fwBbMfQgIsWj11o93N811a4A
PjTzDLQ/mlzGtrwkv+GsHEU0phSU9TOtVdRrVQTK7fBlff8WjTaUPeYdD1jwHdH63pbHkl+k6rXl
XbzoEPPe8Pgh01DOs8dZR0fYI+rlhtnfWleu32T+x1KZ92RC+eipEP3oY1szajN/cKy8Qhn6kQFm
oPOPHZ/mepmbcSJ8nz1Aveoe1NCR6Sze4bnv0FW2lMypO9x/8jHUv9eOB+aGU2tIvLvpSLDWZI2b
P3+yCsJcFTIGFkX52RxtQCWRZom3t0/BC7gs6eT5XzVp3pPGFKQ1lc+GuaQx/TMXUA0jdIdcIu1i
GAI464FkJYiivG3Of4t1w6/DIEd0bh93eFC47/g9p1GNONMd11EhrokvaPOPAJKtjwOOhgpUDecp
OQVnObvvxoN+W/GxT4k1uSNufrbhfthzs6HPO3yG9s6lPne1tlMbsj2mT/TswjVDhq0o72NOn+NK
9KqJwjcdrtGPa6FMvld7O3QPzgt7dcRG3yodjU6gwBKLFx2vorbJMOG3kqVN1s59F9CyBVQ5XokW
ndm7+GubE0BKnVYfMNIZGIWSWVrGSrFtH4ZDQy0lvTK9XqCoWrYhWxPmhkDYYQTEKYMjBqUkbuGz
z8dWSajNUWC7B81ciCirr8+VIfcFL9L3lblnVR88Gs4CxFHHfh7btPnFrse2hCIZvcPmE5sV4ydl
jVFLc+dRew2yKUCNcebGHix6bgMJ1/Ub8baGQT/WPCPscGjscfCq6hPJZmPWmk/Jr1I3fZ6NudaO
fuNM9ncMwvKdJ7IRy863Me1VL6SrwEddPW/E/r+GS7C/+wp+8lwqb/SHbJdrY1gYg+ChicX5Ess/
5rN3KjN0dA2sfex9dNzHxv6xiCefv/AG6TJzJWSVhtU+CfLaPQyllQcbrWxNjhFsxE1g+58FKWq3
MKUXYjKkswAdZEqUlQ/kbBtWaCyjr+fbjqG23wrRaRrkep1DthQpVpiU1IGXxgdATXEL8qlGtScM
MopL4HMHru9xoiQeoGBYmseTZJjhGRFzbip77Wd+56vr05rYOkRhui6XwqKJ0X/KRTViJJk2P7T3
47ig/r0HPRyxoJjWGnWF3jwRG7jMFAb3kSgum5j+2fWAGKQSYeu3KDxqFJVf9yP2hCJZ2jqP8Gkr
uNdstC+YNDr71vdl/TXDSfYvcd1DC4NYkITOzzyLHKVHDrLpDiA46hQVXvMVFEC8N6kbwcA8llAi
tMWmZAQEbTy5w71KZuocWeoT49FWskcbubtLsq3qi+GEMyo526in3Gt7ii1lm1dR8h7ssJPuHWIJ
eWovHxTIl4W329NXeu55Di2xnuTsTywhow9a26cQ73ByCUIUAgWl5A536Vrpso5WmCXTYUBpjjF2
oEoP8Qos1NSQqC41o9dsL8ze8Po6+GTThSJYb9p8zZwMizRHEcc0lKZcOIWz7qazhl6Gehu26NjG
saxmAPE5gqk8zAHYNM96wYns8WtG2VwoY2XiTBElLRQiwiloySgHt9L0Kd4LrriJG55X3r6f18Md
TLDlrT72sy74KVKxubOJZhLfLDWcP5AdCK0lagQ23il4iHnDPzjEFaFCR/2gfM4wLmq5wDgIJYh7
eU+uiLGvZBJq86GMK2BuUvM0zWUDllGxYdds/fIIRdkIJgRuroNhifOaCmA8ZGI5VuHx1s3hACWH
bQVn51oppSM/e+27yH4uX+2LfTqzTgXDS9tsotQQy77MmzQoEFV1xexP03oqoJCXbTray1iCIOT4
d/lcG0U6Xes7ZzKLrPbV58Bu2eZ0qtCen/V+ecITOERU/Ap0TMdg/XI2Dg6SH8Uqe4Xq+2B+nObM
c47TulaoEsZkRDfbVDYhTBBLb3R7IPycXf3nUOUYKdOwFOXoC57PUNVS0iCw2n2w+XQ2qMrJTozp
PZFO5tggI9oKoZfQHVUwqQQoaL3Qbk6p5HpwJ2P34rXl4CP3keCD+U0o+lANOd+PlgAowyEXcVWr
+nP1MaU5h+QPyxWWCF9Mjr6Zq/oAFrq7jLUWw/1+2Im9RCi4yOZsrjT8fitf0DTf5GEppnV+tnan
w84KIXdESZpwnJmo+cZ3ldlFCRCizidKq8nupn74LzvsZ/HqQnNk4HzX7lG+GNyd1hNB8rr7SAWt
9Hri+52ngR8tbeoMHnjAsJdgl68zeUO6gfhXKZysBxqOzKa5YER1vm910TQ6j760H5oPAx0VzRHv
TXYeagnpqc1kdTBAxA/hjfLty4XWj+/sZMs2XFHRRpW43OyD/W2XqKcw+PtKgR5Q0qNqLesCZH7a
PT/kzLLILr+Hw7tkR4PfUO9QJq/M2Xot7a0I6JYOI3yx2di55JYJn7KVfej0hkPX4eB+WCVtR0sB
3/z4dBlHeG1iHmX4Jek6RQ2YzMC1kJSJLheMRuiDH7ofoIXy2a6xTH6GRhDGEnPFPRTfUoCIEOIn
8YUAgiJhBK/qlATlQbyVGghPCDZKic3w0ajWDW4bbwshNDyc2+MRbHNXLbdzF7MeVrlwmgLxGQI1
a7sI67GvZknWTpNg23NP/b+GUmB+bNz7Abzzvp44PJ1d+HFITrpRP3QsaQn692vNj/bR4zZdocC2
unaOPs5RzfWzDLYInJlyZMyXbL13vN/rd9dqB+nhUFMeKARgpufpamrS4YmAbX7P/k1AA/NmLqWr
zuWOlCaqVa11XfYEt3zdXXdi+cvXHtVIsJdVcP93yHIQIBhhAESeqew8pHLE57R0xS8b7eYq+5Lu
/FkK4KFc6WjwmXjHxYRmK92Hxuz/Re5xwNEMWveHQu+lWReHQXhPeeK7MN+BRkE0FmTR4sdmrlci
Q8hrLdg75WdrEOcJWz5xtRMpM/vuZuoH1L2Ndbwn1aiACWI8xkbQee2ophytb4Rgf/4OjLSPDU3B
s+Fpa79UrwkJf2LwwDpg72Lu2OHgqHKk7WCjwYRsrszdVJZtqBHaufNRPPyKleexM17InV935chF
cm8K+wvzkKoyAWz6n1Vklk0QABV8vp3e87YgstHwVtPoPUQnFBHFthYngxxubgFMlzby41v0Bmnp
SJo+PcbwUjbF0Ser/ZUZ8KYCaT1TK/qpgTGYLGfC+2kx4jwLg6ZikSSUMKfybP7hX8f2OqiPb5eu
djQRb269hZinltGb3iJHhX4VXzmv+7KgCjb+At03qR+0H+bHiy7wI+dP2XyMlVdrYFIQK4na1jsX
tnD8BIB7j992FENo1YQh4JYkfRDjGdyWYVY25dXlKlyBeGzl8TDGqdW5SCXO8l0Zj5Fdcw+AVe/p
fQGTq2+cOZJBvpbLSvB3EVn7JWVKwqIPyA0GMD/z17l+EDJQ6iwROSUWtvFCLSPLERD7/JvAiFe7
nQ3LCyEqZZalCylRDypUm7LwqQF8bf9XRkdu7bplWmIEirPMwUjGMBh9I8WoHx0F8bVEnbcBxolX
hIS6Zea0NXp0b7pRhA2/PMp6aBFr/yiLfX3LHzCN1MRVaoE5CWztSd2dKLUCqLVqopyro3jDP+Zk
uod1Wmg/i6kk6QDTWkEsKuSLKzHsNm1sltv+mcUZXBpXxYdJB42rK1PsFCUVcdOkKcQeK0LBCa33
+BbD05oaN3Ax5Iwk8MeFIje75E5mo7eoSxLDH6I0bPV1/eIojMoZAL0Y73lyYm03LUTU6IwFuW0e
zM+A9NbV/5ALEVmUAAcYcMMfOrxyIHI+XB41SZlkNAtRlsy8xs3KZwHSy7iB3B+yw61Lf/mIZ30V
P1dHBV/beksNWNknyIsZfYtDBzyVN8KciF5XJKMvK0rg60qKPN7jHx5dNXgPnkB67vAlrDV0/slx
wHmr606Ah55MHjPiQgH8vqroP4I5rf1HTG+fi/rd4h+7x2RrSkh+Hu2GhkLEEYB/t4sCyxRhSunb
WDeg62oCxfzpydbx6MSNvSp6Ofyt5qY+AojvjfgR9ox2Wl+HQ34TaSvj1iLHzNxO/xVPtkst54DX
8Z+ych6Wa7VdQXdRTmumEGE/RNbWOinFxKMMhJYD6UBCWN1Gg3hW5NW2sRbe3O5xAPEkgWKofaU6
eOrqfC8w9rIi6tjHZfzU1BhPvFucPLr+KLx1uaaEaxW935BAyJmTnJJvXdGHjnRk/wNrI2xCpPSE
Cy/6dtqawePi3bwsVYx2w5s7WlOBK51Qhs5a7WsVbA53rl534uTTBeL7QYzpqv4rtyY2nLdn/hZJ
r/hJB8cw566CADoITdTHM5MdakMU7qUQq9MY1eMyA3JncyXfgpTW7xzagJ+bPBFhoJlb7jsgMvCm
mgyKfRiJecTxhKZaDUb3u76/03/JSR8YjIlnQ+ugDngakBJ0D0+5Jy/DmDYhBjV1tCjMKsjQl4zW
5PqZqk6JSH8QU4n/G2wSABR6CMfWZgq83WhpkxEcL0tV3zuwxL9nRS4r9T8ur8uLBk0xVq84SUM4
uvFBBYGx6lvcJGfN68fSAfoSge4MN/a382QSltYuF6ASHi0E0S9jECPUpbwG41KQ0x0Vej1c4QDQ
240pkHj3OGd1OH49oCTJDoSbeAaQTDCy9Tn8QLtaH6xPoLuRi0exeU5Ep6RWEotkVIrrzX7zs/wp
0bx9ilo+hVGV0XuBzKghz6iBvTSsUFqMDXQNGLzksrtpSlXWZ4crSzkrj7b9IBK6uhKkE/Ivubny
uzkrJKbhsR0m7jdkGrkCDo1AqiM6qhatj7c2tEQAEvOqDUqqL8ZYYmKvemF2ra6L2w7nU53TJxs9
nLfhxbUAj42F3DEfsno+eRKZokibH7FIFYv1OH0jh0xA+6f4GcDC/o47N8kWZIyUBfzC1KfwzMmS
bzhI0cAfS6NjhC/1OOMwzr+9ppBMoukH4HMp3Q0tUoKWtAAd5a5HksOBcd0gZW+hoGhttnfTR1lq
b/Pc440DOxav72URz9ZsK/sRrkm5T5DT6tZMXJFDadeDenir1rfJPwFUzya0RDqCd+IotlbdwYz4
dtFsEKVhM1V4xCxXuywboTfBmgFHqAo+XRcRoLzqrVYpaALXMDYmKadBl4c6eKSOvAuHZsEnlStX
9jaCVbaS9qbtsjN1I6d+COIWhEC4zyfQtDF1TgpkbtptOPTyxfzWLH1K4e1SZzlkLvxpLoi87z+z
lEgp4zLAzVuqGgeBo0NwLfTb/ZrOe8tWma92YApXDuPXJyG6cBnqlS44K2IR6NcgCz30+1Ci7MQq
eInaRPtV2xmM3pQnUoJtAJwRs9JTivrOZwb92d2Rc4/yKfWxhPw8M3wyGVdvc41B3PoncJ10tai6
GToDmMl2ziUDCpBY0kkRhLdVqz0taD5OKvD27R6OsBRQoB/6nEGqZU2fRT6Dc0Ua+qp6YjN8R5qy
ow8criNVKSssQGxegSyeqVpPvMiHerNf5I75bASvbDDU7e4Ole4Y60gYvSMOcqqgOiKJjHbmwWhZ
rVGyaiiKFpTEo7P+qaz0TNRK6BOXRmTXubGMf4/Yih3KuD6Dsss6FvUggwMc4b4DYnDop5y4e7pV
cux+a14bEwWs/JWCjDwFu3GtpPqfazM05TNbEXM93ZaCGVAov+oV8CXwu96WU9nzaOGld93mTwqW
6dcpZ7x1AaMokzrz87+r8am5rfT2TUwH7fCqjPz89E0hGx9MwDZ/p8jaT90cmwSe6S/5bi/zq5As
4K80ep7s2Y7dT76yyQwdLXR2Gyfv5v/oUbt6nc1rpxvpZ3XFJni1EXYEFaz/2F8Ezphk4egI1sZG
KLu5EwWvV/oxlw+IqkZc7eFcIuKo5nFwbrLIcMgOktwGySb257D6KXDYhiFIRAMDHyyBrE5p3GMi
yrXEL9zTa2qR5bj9m0mlKJnFuutf/cFx6Wn4QrIva7dINnJTHuyw7Rj13lzwpCEVaZUh4BY5Ysyy
F6/Qh4UyKgX6MBB73gArnsIr7ZzHgMk9fWVrztty8HL+50hppgW2MrSioa6VApJ4Zn+xfkJwF/Tq
IHxXzSO5XC6AgUrHOzg9cyCibVmPuu+JIDJprnspTeUVNbd7hufhZ2v/AkWKL2C8lSfNFkmKx2fT
xxsSiSqpyA2cbd/3wnFH8LLINNMALomKVxWT+8WOSS6SCu7KBWc5DBNCTZDrVBA5FPL0z8gIw7dY
XMfu6Fo8Zc0hZsWx+IhaTzKZ/O/dxcGUI00TCWyBqWZbedaqnYgQjgM07cubTtjInMmf5UkBVR5+
H0nnCFt1/9JTFzlLEX+BaWgImgNVHcFcTWcJB6mw/iu9424NnZTgUtE/mC+EDWGFDeV3MiBVYTGE
mHt2cVlRM4NWKJgSTODPvyKfupL2SGYQR9Wo3o1izuPmsQCBKUJDc1eyG+wVz2NuGZaef7qCJ6rp
5alac1gq1sQatfs6SGhfukEstz1kC5yXyjIQb9XlE/kvNLykmryTrmE5jbOskelGi4UJ8klWrkUF
OSbP8VZvcUU6kZglf9iohsUWZm80kcpwSahn1N6GQF4qNC/A31IGgG43J4XB7/sXx3oxXGW4HdUJ
FM5XnIg/p5kS9KUrhWwW1I9qzoFtnR/FQ2/5z8RKQ/MJa83HRWSQNbTTCN/Cz7gPucSSGP8W7WAV
WmCXirwfNqDSUNZhpMOmwujiqjWoqBp5XJXVZmuxpFt0AtdqbZwIJOAuTNn9KoD2nN+TQRZdazaR
ITrGq3HXN6maUEMtA/YPp7yc4KEhgw2DbjzMxJWPYJijyErqM+kCLJf83cdRWP5IvsPp6TkoRia0
IB0a9PfF2CoixYVJ6QaplqcyOCBDRdOTgYR0nxukr29L8doU7nHi+GNIK0QKaAL2x8qzC+zo8fA5
fC8Bh9cni5bTd/yAmRkYjLFRobCRWjAYmaxg6hvU2yywTjd1szJBssn+JdwVqPfWuP5g2tO3EEvD
m6W1bZLgi1NBrDrzDl8dxH7DqgfuePwx8GDbEA4wIc8iqjygWU7mC2lFpJOKDJZ1yI5Y31eY86my
LqgtSjFlygC+KIrmXx1MdOPxeWmQiaXpgzkY2TRKV3BXY2jtwtkSfUZ5qRuNUtweEEqpze95q/yE
QRMg2BH7tWchFOYDPuS1bNTEdOXQFDKymGztaekjmXT0h6n+9oMW0NzDodtCHSCy0a2ogPRRFba9
qx6jtUd5OJ+HLsuXuwRFggdAPMnRyAJG+WfF3y12ffhFbQCSGR9s37XAAIW7hWdH8YIZK7R2BX6T
oIlST+kxb4aO5j4+yXjcG5nNkSlyZ5XbF/sGPTXpYWPjgtoGYct6Wjzf/GJ4J0jpA3qKny64UObW
dyW18rfBHOOcpmSQH/OMh5gwvJf681EKt0p18oeqQc0u0f9wn/0patjXdXQI9qiqXiFoXKq5jxmu
KEOItr9QXFzs3p1xXwNBQ/4id5NvIJLdBFO/9q+2HQINpqUsxN/DhKwd2rnvyHKbTn9/pbCVm7+7
9i0Oj+ubzPOAxzHJKV9pV/r/X4/3GqgkAUo4JySBXvzk6h7xJXNeOxF3NhMa4nTZ04lmMSsoPOp7
TVG8nftJ9lacZsDU0VuP0YxBjOmHM+KuJtFUlajJdLLazKPeUIWXjMvb3Uuci2pMROOfItyusLdC
RVNINM4O9glCdVguYFQAxhqXdlb6XVZYgkhms+s0mRRtAO66tCBR3RV0jRsrqmsoWYIhp4JLX6V+
2UW3NFfYSsnlideTttmJpdU96TmEFT3JtvbB1+sVlopYwgMNq4WpwC+v5CW43XCYoZSAFKJs6j9N
9TUIvrxyi9ZEHFLbGrXon2oYAikoQ2EEkB2cleq+5Hbtdq3I0Sj+bLGqasF2iISRTbJUykDLocLE
i9C3MIJOB4331ORLd6gEq1CogoMpPxTTCx5pSEsvTjIp/eUuRjdWJloElFj2oVK/8Bh5k86UoQ1I
FtoBdSljY2mVdowcCLXw2y4Dwit8nmeMqkKJerQilbXMvHTA+be+Hm3zlR8vnrIWV5gVCn9PLzfv
fQWdyg2Eov1mJUwmv3y8kZjA/I+G5zz3+0lXuyzpVNqG60ONIHKpxQ4M6CSpNYGOPQgnhQa+Q6m2
IE9YsTgrNjGQ/sV2CTwNir3xzfMi75Ali/Q8zS6MyhzSvf8kspGyNFcErBgwFbEEqY0a4D2ZFav+
jKNUkydmyQVOkt4br5vHfvokQ8cL4LHg7GZc0SoW9nwLjI+JAiVe/qaqWenyPw+XUqnSKVwPqa2R
+9EF7gkzKLTHB+pk3UHicEGGaLXn1ZtLsN97GzSaGhxilQcJqItCDCc7G7OJBBZ2EYB36NLF+HK6
AB7bd8YKIaqyYNCHaF06CGKogOYWeqd/jBlhgwDbSA/mlurBtTp9rYs70eVq7bdl4Pybq1Af63nx
Dwgg0pkvrHAZJ4FukJALoJLA64VgQ32NB2BA0pvuACnfaON6KxuwKuyarOHnt+wFVc4jMjOobUmr
Oih7jMEOuSdeLHFwFUtdbrwTtEIXeMY++6gVOdvX6pqBLt10G1/eqnEJ3NmOlp5QWBqYUNZkPcHW
VDWCZN2jHLs88FGwg2Mne658WRN8NkhzgCueENUngpXP+6+P6gZzvAfg/c5fva5Rqi6jN/5lT9tZ
wYxCj/EeYztis84hUTcFPpGg/PrKW6SpPeYCgHGB/hkpH2g1h+IhbKGgxjM3kJdDdLkdokEJYqjV
J1AWpDMgRHuDeOAHiKH0qsJvo8kglzM/CTZkQulkfdylJtAWRfKlWceaDGt/d/6m7tBUdZi/ScQF
Sh3fnd58n9DKhLlERRR1Ov0KQc16201Ps3wotrkRuFX7/KcSpcHL0XAgpz1mKrbLPUgOYZQGT11x
QbJkMOB4hCL4WbsWQOWx+ndrhopTLB333nf0zg94bY8y6EoRnmaRRQDtF4U//jU/3vLwhjX2ls7F
LQmqXgE3deu6EgTDtpwWom1DocpJQ78isBey8xR5Z/UzvbXeM49pwAJfXqAK4XorI4m1+Vuj1xIn
30SqrvwoTHMmg4W/NqIGVR98rlP2YDN7/izdcL8J9bQqxW+WLQKrIt+IcldtkXAgCDUu85xe+i4a
yXWi6tYaSakLK9GQzvLs/9A7cB/n0yQVbHDEdWNBfZSMZpWgcPuACwoUSXbnXUhyNryK4YgpcfuX
5yjtDzsQKObHPJiKYp5wmeeP51z7LrJFZhifhXdaRADCtMb61JxcXDj8rhVheiYoq5kVKnEBrZlt
FlXjRc129lNL+YgO+WiNxrepauhtdr6Z88Xam27Q0qWaA2YISntwPSsLN3CXUbGctdew7CHAN6UT
z8ax4Ynv4IJY6dmD4BDH+ZEfnY9XZWd40vlVLeOByJg/PsyNmAwJ2vLeSYhIvI85VWBkfwn9DOl9
DTpyWcwHTjccN0QW/P1iwSQoc4aagOFmoy+1NW2EHscbbgr1eIxWipZTZXjH20Og0W7WAYUGti7o
KKuQ5SwPDkwA3UfRpnguOpSmmgdYY4Iu7cXBDbmypuBwhNbOCEWycSqCK2YkSQMwqIoGWBcUcoN/
vNpzzrTkvs/6aVQbH/La+nxpU8L4RQ9MvzG5/zd9Dh64/Q7D1MY0/eupubsDO2FK6KMLaMlS1xoq
NTzaPZRt8NU4PPCptkcwiqNeka5Ib5b2s+o+fSSReXHM3hp9/cZJchE5c2yDRDsw88cu/f/2KQ4P
0seiya5K6IrVZ1i+/0uJMUaLto7nvtZqgBiqHwk4iuKXvVPI3kJTrQbEDPR2iMEFFn5AoFa3vqGR
K8nghtvyPFDBwjah5rj33JoT8aeLYO4MYHcUSVuMaaZfxsUUIRGaG+HQHiJNWgO4wIU2sM3iP6CW
WIFPNwPt3DrOnmOjjkQPANE2yoA23MMNzDlSY+lTUVNOEGDYCEHDIQG7zQ585taTvRzlU94r+k/M
AEIESTN+tqZSAI/AdLmm06nBbdmfGEAdBv76zsEQHJwCaPeLpByXj24/83HC4dnoZLMn4Me2EgZ7
nm3s8cCnnFV+R2PZrakgj7RN6QPuUs+K8TsxHvDuW0dIoYDPMHBV4xiUmsPFYUDMKkJf+u7bJPal
N/pxpGS5UQA5buAcIRLo4fTscHphXW2Kam5j169Fzit6g3bVCFlj7o/3q8+DUQ3xFcsRpvDG0OhO
QAquyTRMg0c0yAs+Zo10iJ8h8MUmc/vlkcay0Z1xwtCS1wZmCVGm4EEvX3VAvM1wt1g8xKQkpehI
6ewsxs8anXUEPsMBsgzNiG/FtQjYwaJUTlGrGe/tukyxmPPhwi/BYCKZq/yh858SVORpUl8ozJgn
+rX2KeX+wtZ03OsH1+vLGrKQdY9xgAkvnG0agipAKU6GUS2pbhHeF4/RtBJy4xovCCDbcx8nSD0k
uY4xf7CGi+Hziv0kphImaIsCdELAWgKmQLtjNaVFhQq0Imuk/opKfDx11NfaEaJHAuM58d3ACE+J
k4d1osvXTh2ITcYLYoWrmL9zMS7HeMG14apABNeB0PyI30W7UwdQNMjapd5AejucuTrggRtBgh8u
3/v+EQ/PKi5UPU7jmZsJnTEEIWlJKa71zkxrXzUlN0HVAGgjjzfDU2+WFHkWP5xVFZoZqlCIZV4B
7TkXEdVDZ2A7P+wJb/tJM7sqoK1Sk5T/RoyUmx/FNMw/FRSCIW7CzScCu28VJJC0b0J9o9hwepjh
GB4162HB7WHAKdmjzHRLvo5nIn3pXOFnlvaCpbG1N2865i85EvGxGmdniAuLqkiCD1KP/DiFiDkV
uu7u/RbqXBSNeXNvvhcFx5EXzaG8+l/1PTcJiz/QSSGF8gt7yNaFdzjz7NaZDtVFvtaDCHzVxHBq
Sm3eXebZLmeuD7e3Z/BZNM90DRLozdK2D6PYvVZgfOdUwcoWBBJ+I93MJBQcFbVzpusSTxlnbN6v
CLkLdvgro+O0QMQUgYemzlYF0WqLhzbgoG/CzjN3eca2pgD8CfYx0e5PNr4O8d7AgK6JQJyfklX2
+E4HQCW8OzxQ4Y/Mo56ZHd8Jel2XJPU3YBRIQ3us6U6cxU5Dwr4DUGkDrHwoGQDJblxPB1n2qCe5
vRiX6C+CAFAfRL71gfdNGjnEDl05NcYTC3RROLclDhhPXYqscD/kcJ1CdYjibsZc+HNmn4UDCT87
zw9z+rT6qTa8l6QG7WE66ySfnY2btZYeAilYJwdlE1CYMkxM4dNimP/RkMjFcOyDzWoTEOC7LdKm
wdi5zpAuY+R7c95Vmg9ZYUDIyRgO8X6RWKT+4wRtZlFfjcfLS5GTjbIb5JhzPkfB7TAg+QKuaQrN
a40d9Pd2/OGqq13MuVt/EM1uVBwA2JR805cG/AUxiCODz1LftJjzpvSwKzJxSWCnTcOaPnIiJ2Gs
dI0zCgpH1EYkXeK86XT7pHV6f4ZRgRB0R1x58u22+9UCCTtR4IS48PCUHztvI+vAUpHqrh1X5vYY
gy5XvpHKMZj8oXaCec7DV/iVxZ+aQi6M2Xm3Um/mEyy29dIaTWuDnP5ZkB9OJw2Hdk3lIJY5Du/w
mp66K6cPgN4F0a1kSYYrb7b9WfH80NGgO7Sq6sSLJmtiyjmBU7PHfFlQb8xqO4bg1aSTwIMjDR2r
HoKzJq3YxhnZmTOpGMtyrF3rMAiUt1prAfLIRP0ZjUVlGOV2DmKRGEjF0KYiZr+/f3ofj6AMhLaR
GrgtLtgoQXihiWYedyqw4L1YQZTEy/LXe2aExG0VqqiQeghheTpKZgZo+c6+AA97sqGW7/w4nzBW
ITfB3FPRU64ObfxhPe0OuVK3lna+F1BUesPGAoQkI+OggX7zfMduXUru9aSsgzBVGw0ft9LDoVYi
RKAYQRvyjMUy4DqcDmB18tMT87Hx6Bx2xfsh6IET8roMWpnkIhoShC+rv9D/+nqmiiYgutHK90t4
zdXduwa3apLdvweslYxtT2WBjIxdKOmztYDof5hOcYUAUuriyPQ+TZUw1nxQsdiUXJvaVBUulW14
0ydHjp9qUruCjPUv/PfNeeu9DzSnw3cwC4CM52pu6O2FsK3ib/+kqr0YktCT5k6XGTjTMaCnCqHc
vNR5vLL/q1UcvTlls0+ET+PPJjkU3veblrEOYc73O4RgUwJ2kMP4CAIAtIgevyFAF9URMEUhp4lm
3YIMug7aCwVx66v74Xe9CIGObE6httx2HY1h216J1P5G3kETyivssIqfDw5gdc8rUeQs1wJ/CAu0
/oDR0uFqRaBUVXGG1GV0eyDpXEwgi6BWyg4gPH4kSnXOFrzLRyfKkfpOKcem4fWi8BzOf1uUib5M
ytHPio/uWm8XeouwyNZ9sToq6laQZBIDdwdjzNMgiAIeC2+pYTpCDqx23AXsOrmvyxwy2/EcD7DI
uufkCXsijIbZcyzVUE+tDS+WC05Fqr9EVE/zsQVZN9zOioIFl7QErn8ei6pUN6P/hJ1qpTkN1jiN
/uFh8kHkXTPuLfexNPqNdDFIl38Z6FgxHSK7NcVJTOINv27q3MJH43+rewe8z9ziA8naf3ECVg5u
3yptg+3Ya0uzTtuHzElkXhN9qTzofiex1/6hQTeFh8sO1rABRbDFoQc78O35Ajko0mXW5fVLVXZv
6l56C/oj9g38kcJTXV2D+7Z5ITqNiRHwm9RbMWNE9YmN9KE1Ax8rXNWJR4HQpUxuTP/QzTJm8ESB
HGWD9u+XGqTRTC+iwYgPkJtc8/nOgDFiZJhjLDOD6KY4sl2zsFIV1Wqwo7O1/UqgSGVba3MkInJz
dLhRewZS/7D496fmy/8E0Uw/XGVqwzfaVUE7o2ZuC6oTOJlnNjqePRBFt0MIbTEEf8F/NGzPxIQ4
3+FEuM/UgmD6NpmdOr+KLP+G7yM1Sm7g1DLtveyAB6hKy0VoQXrlkXXaaLn77mHazhB4bkdOL/F4
40AwD/VfufAEDuDoVir6jNromgE/BL024WJ+Vx7whlgrVCUWj46d5JxTP1mQxysj7N2/IGgMpicG
0Tio3XnXyEXA6MvqCxuG0ELAsG4hkrNrZ/XMIzm/uD5vYEFdOa/rn9AvSPhYTlGpjC/J78McKpL3
TKV4fYampu1W5cLF4bzwAaUsUp6hvIOu/jWHlkBsorqMWINiCxYZEzdFgqXo0MbzH7YsXBBeDH1x
PYopU9IY87VfyW/OJBXOKMODSMMQ7ZbvP72IW8DoQV+RJCFDf49tEZeiFnfBDGjGrk9fvUKMw4Gq
2ocCNVQnDzOFIjVktGzZQtC0bD8UIWGQltaqvHf58LfzGh20O66UszM2CWoqJTVEdIRUEp6MR77M
Ri9Fjw07ICbx0oQjJ5GtUyEjyebx4gw1kejX5lVa+TRicyJCCKeagGAt645psDCFpyfdO1wLBWpn
tgJNRSPo//3WiEmVBKvwbZYFInu/8jdPTAqaGh7W/djxukGwclz9/h1Ba4jDIY1wrV5mMv2Sna06
5vR5935VHRAcUQ3Y4y/0bgvHR00SXMlOVtlCS353aGQkDm3J2+EkMClXJFNMsvTmy4Me8L7HFvSj
lklXA8OJFC+5g4Pp/jOjlKPtNmPuGcr/F+70DmfyxYA+Eh0Ug0LXpGdeUz2AetYIEmVkORW0ZI6O
4a24g9kiie68jghmK42367wuiP0Qtk9jsu+XSq6SBb5c+rFyjXNjpRdqLMsDwo5uiEwDyTFhGhjo
Qk3IakO41QziLjF8QNaS54BMx6ETW5TzvyhERcwKykYH8FVtgDCpyS+oiFIJOSdmZhWhpz+bq+cG
ilG6y4Wr9X96AU6fKV2DIV+t0fjMjcWtRp/QXo2iGw6Qj8hAw+XApzTmcn4/2TimU1Ubydz2pzd1
7B5woD9BGP+BSGBVwmOJe5YewHY7MYGdEq6AV853DZQxhM8MWyNm79q9Rt4uudwsd8YJ5gGiF6wz
ej830nfyRpOrtBBXwXiBnQLfqd+gOnk7GqCQl/IOwoPWFS82mIPR52Dd+eidWHwTAG5BoUzDaLzH
nDMzkJ7egFowOScW77gUCVSJZq0XdnfOTHsX5dRlJfOUWQByWSWGPYlJ9nYke7s2nXZCiIU1a5tL
y2VVXqkGq3Mjo/ToCHT8VFQQsbiV7D6IQckralUIEQIhdRz6MVKEZRxB1n2BhgPNf27LVZWwpphX
UnM7YxfzpLkEqoYlFEUe9jh5539mgyrXnsuZBxtHjRaMFxL5kl9GW+TLrORomMP9Ov+ZLY+MwaM3
SXMGV5F3B/OBmc5K9hd/Qt9YDA1Q4/i/LwXD15fERbTS+dly/98u6jOtp8wwCZtM31Ghw27rnQir
eYUmGOqSidDgIkX1+4ks4qrcPmF4mJ/UOcOGXMNmNG/eu/nIjaDPJ1ZHx54BgZteL0sbHk5CSs2O
AIH5WXvqGXqSQ0O5rqrOLcXM80Mxet6KAOZUTHQYdd0tKpyJG4L4TYZqgmQqbCs8XuOImo+LVh7R
EoQ4iOQo9auJXfGpqsH0TgvCmMUsdTeyzkknKpuQcgsMSTDQ/A7vdzAAZr4CSXeh8ptgxJH7NZEi
q4N+wut2Xq8+uFdIWl57jmPuZZEMpGx1CraoHktSaOw+nslzn4qPGVy+Zt5hSfdx2UpKOt9XI37T
ynhS+luWdtGZl7GfeqxobfayrKMZdaym4gBhxNkN0mxpu9Vy2T8H/cuqbAY+ChERJOdw4RXLI3kE
sOiRQCNaitsocv28LGl0zZRJrNN9as6366IpOnqIRz6dV+S/bMH3PEQTQkUI0aPOrSGFRLrRxxoV
WC+HamulsChjMHqPYEYHEETefiuO5xtu5Er2l1rxTSG+h2P5iD2VYW7p3s+FV0H1fw9j+xC/x8UQ
wDiqJ3lGLK1Cqf8usUWxHK0buvWLq+Y+6QCL2ZENc09KN7OZIr1GRm5P4pffJX+CZsIiB/Mbln0H
F/UcnGyDRXaQ1rDt6+It8q31Gj3Ptp82uRyQfO8jRwlVQJZzrI7boKoe32E/2Dd50Ca/4sergd5R
XhApI9FKw9/KWblsPvMTx/R6GpeBYRJLvOxF74ey5DTUByrh3SEEOHRsHuHJbHg5rNIzqCNUnd3r
Q8r65K9+PwWyguf4ayiuT102ZEjU9d5z9K2VdfJELZkteBCv0/IWC4kcF12v4yKI72zZBk4DKH33
SgjISSdZPqqrakInVvZ5qDguZwRYOokOh0JhOf59sVomZu4sGXX3AN1TnddQa7xpG0lDfJlAEiyX
I4qdNmqBZfUW1kqgCb6V7bTRn4WcxuiU2GhAMClUJePojMhFBe7+M1GHoQEh1iD4OfqvpbnrNgaG
41SY8d6muCa+vW2XrGZV/QVbcZmx7ugznxnv1BMkTdfAMpdby822BIKWIfF5Kp9CGkC5PPXyQ4Fd
2mMqoNi7/mxM17m7Kg2CPTMWmLnpLGm6gCe0UPds5hT57KJPlZMEvM5+iCIFIupfOc76HDNP8Ixk
49biSkG++oaY5c/EBcrgMfShdciFRh/5KIlFe+yixd4FfHaBi6sjYVmg5SstxeNIf8ysMPVpQPSB
gb+G2dFHlqPnrwZ8M5Zp6e91l3BOa48Lt5R5LsDaf3x8J5nKMHE6bnoPggsQyVPkXgI/+FI0Vhll
WXB31M9kczf/zuXsxWSyQs/A1BuMf5SC+PaBpLrKqlWSg0jYIB83bd/pr6T+XA/J/WxOZT5p6B4l
8PQtXuSCp0wME9PKQ8yknGs2ay341VnShUXrWma+YzE3gqu18ENCHF0vqktubvr/KdetGA2tkXiV
AF4Rz/eIMt42nwJGe8KVdQO8aMn3nlFY/HVcWtHUAsVGGozHq+o8jAR0Dt+JT2EBhl7uMapTFmoa
76oDk+BNAyAOnnr3wu6hg10xXRCPnn7sUznX8lDeAaKcGmMguMMjfl8ss5KzIyOz2weMFZhKNQ1c
E1E8R8d14h6X63qOsZYlZMaZfb1KLZ/c13Vhh2EFsNCxP5zrWYHleesTvft84Lco5CJ+r0SCR5E4
m4w0hv0GRAGSaq3SNpbh7uMkjTJL1TQx+SDi0dVtyJJHfE3gqgGmdFPLlOATgkSZZ05YuGRwQ4sy
7vNn69iJ76TkxtaJujh9wDn/hTeM1ulME1SUSaz7n0K9FovjPi6qyGHabGvLmZ2Yiv75bWJKLaiO
LembE7duP5Es0bSLxw/UBLecP4q8ArnUvDW7W33Jh6mpkf0BkCBaWOyaRn3JNbWFnE684ugmiEMs
BqIA6S2+e7zRmYuGLrAEZVLLJ0Vs+DIaPyYIazO+OFmMmxtfJDsDW+8I4GajT51nA3x6Z85X9tjy
33AZhiWQ/1qMUy5Mc31D+smApb20KLAX6bkbnZeGKZN2qGWCLnuWTxKIhcrqyO1c+ahqGsFy0G48
U3mKFms4TpdS67Ps7DJAcT9BzzlUVzFmN/99EtjXRNuqMJzacPBuHEOvpZkHiLNn9WWz4WvD3dvi
tc0KLboSGEUv7//LawnEjzxNFXt8sJGNyRNJsi2UWCPauIdrI1dWK2+S4GB3istI0hUnnl/qoGYH
WdaJdjBtNN5syHOSPcFKkbEN/mhgQOcK2PDM+sym7C4gTzwoNvSsywN9rKAeSDRMhB4W1ms8WTZK
N679CLbt+s2X6bdW1javN0hMN+A2H5SkZ92jMWR0eEEVMvT2igNq6oz55aDQ1cbVZxu6vA/UiF5U
DBiw3DAo41Abs9q7i4JnO7FFLXnClhCSKnAC8hGBrDmZdRRNtYePFyPcxL/E9AQoowk02g937BNh
W64X0BstycWRSpraTfp4H5Olz1fg3D83p1bIbTb39YCZhDkpgYfPpFrSuJCZI2LNeTJToWkif2Y8
ZXEXRXIyo3+3EoCabdxNalA0mVHBoVhUlLApdWyDFUtHe9kKUSaJl8+ev4RsWoi8rmVag2WDs3Hi
kJa+/Cmctigv8ZSOnndhGhNU7jheys6CAeBPynJ17wrx8xD96sC8aj7LuiO9o5a207RjfeFASNY4
KD2tRmE3gYiAnYD6vii2ghJ1o4sXNHd7zNw5rGOs5PUOJiXbqgnxNSGH1953htsCfoBLZNcDT1Js
S3m6mYLtODifhzuo+9WwNxCZvCDPJH2cyx4D3Hg1D+NEDqyw+Gzw6K74eRyvj3UR1oYSmNVQnu0N
N6IwsKOJ8amVdDMTw0EjV02dQS4Yz6JAbPX/2/CB0HpEANfcHRDNkNlq0hWlQjq5AQ+Bjzyr001Q
cfuQENcBZSLvIuaW8oDnSDj9LSaocQ+Sk17ZccI0bDqcbFyzUETscwZBXf8IQqacxwD8+UXHXlmp
PLI6ZP2Jqz9xVmYva13A79tnx04+zuMUHxss6fcv/izexl1Y23smHlpppnYl9eZw+unyHlh9Nety
lzjhpFmaJ9ppHw62lL09FEoiEAaXCEGpaFtajUhidwduG8YyoCxgnSLgemagic3N4I1NVCyrRBNn
ZCqGKFAIyIqIXSV1QNG7t/kQ6VFDQftPADt5Lxvdp7jNUfEQtwgvU9FTyzFDOj5lpZusyTaGPR5Z
sgn0Snq6CC8EVhHBkp68V/hlxoo/RXeva0vwM1Q9nLe/cUt9QorN41cpxRp53sUmQF5LjT4DQcX/
B2LVnQLeQiJ28pT0jhNl797+WQAz+zM5+pwRbRYjXozY/7AsbDSrqTF+Iox5npUZg5xt6ENY+p31
aMPN9iqytMUQoabeCNaBgPJdDzy7gReR4XyfqhdFVF/jVn1cGqIyv+62b5qN7Huy3LkIHwpPvJ8M
ssC/3DzqTsgBBSwqrDSh/h6FvrAkHFv95paTXmhyvsV9gzJJjDETmW7UkL03bq5N7vRJgPT8dztj
DekSNnYhUkMQ50ttDhh9WrYdEFE56t2UC0cwpYJ9y8x1cLaxaGVDv223UUcSMwkXAENWHMdfoAAP
Lq3rsbnlEVw+yqACz7BnDOFRWNlnLESvA2NGu6bh+aiG1Ja9tTq5wKBFcSLPqZZS01cmXnpiAUYV
53NaGm59ThSjx1OlFcV45IavuhlIsy8VZbxlRhWOfDzD+Nz8jNRDDJBy2mco9CX/1WhAf23W6yza
nNF9DAJyZX5K095/WCUhj7Yz43KJvysOGpzEyUX1Q8BjB2K7BxB9P4tZnMQ8MEfu4yXdvq+4AsIB
WTFFe51q9zJxqCmsd7LfWkbV7pOB9bZAOSAOQOoMAPkqCEbStZ09o2Y0Kb7B5QIXijpr68WXcIVV
HkHMu2NkGNZHujxmNcXmlApCxmFQaf/UE26lT/ycDWnaLyZifT6InYss8k/iuCm43xmiDHpCEAfk
yYyfoWEBeR4OhLF8Fd+yHceAJzdtjECdp2v4L3030IKukkuoVD5+RVjnPAzaLKyTb5p/a/HyDISG
SPDAVgsL3Xxax3eWDBn901BlgLTWxHFGBkuVEYnzEVAreXNDCB8ZjJqRkoAWB+ttNdrdMoGNB+lM
RQfqm3x6APJDULVkOQtaObCLy6mOeyvEER7wKvpfHwVtSSDLusZtzaBUDxwhDEJhM1jvyS9Quqru
gH0zpfv/q6UOshAUy28PUDdsJjHxgv2OSKG2y4WxAWNeRqZOXnOh93UDXXr3IKXuzwV8Y2133qux
eKlKQ4/yq+rLiuSplaAGStiRNf63oAZdmAWAVtJilCAWcq9MHLhrWsQ+Gpf94mJsU5yxX3t8AQFF
DT13IxZCrCxCez4VaDPWeQAsmv4BzcCByNgAJuK6fn7WoB5qUiCwl0Wtwn3XQf+xdsY04AHDGsoh
sRX3LQPBH61gG2DS5AEFChb9MeqiWdSuS6lbMlQqkXzKyxUZlK0FwyLmEhhEu3/mqj+ZgF+DIzWN
1fmYi1fk3iTo3tx3TSckifF+GKWcnQNT2LSrSYdvM5wCZLODMSP1TKPVajk1Y9A5dLXpy2yL8mgF
1J0NmoquqzxSVcYwblP02YRWuwDOwXQl5UmPz3+jgZSSazzqASFqTaNryCRkaDmhUiIsh7fNOiPK
cdqR2OS0BBt+ZiOo5WoRv40tZ2ofOo1FWIUoM11xr0U/mtu94DgsvbtxuJGeHveRt8Hq76emw6r2
1sm4h0bG8ogBqAStqRdKRs29Bpan7iAqL1At+a2VX3iPd+vg0jG9YHE1IRhQZNsZPnaTqinfkzaP
Ui+PJwn9igJoTjnj7LymFQ0vJ1mCuIbrcip/NTQpFm6r6nzDwfv1loDfpLnM99WcvtKtWd33tavk
VkUmtsUWPxa8OKHMUf9575pZwUoxzNKHV8PsU8FT0yXBIJZ+QK20q9TwGeuT5LnI7dXGcmeJiMLu
0CkcXWBWjAJG2jfQ5StQlGUvNh4NJSIT56gESEQt2ClzFCl46j4D3Yb06xXxi2OCrhcUfbmTeAdX
flypFla67ftl47pPi5tGiU6UNi25x6A2iCmi7/xCRx0JMINQbWbvbHIdHRAK+5RXsKhqNsB2jzN9
gbbOhr7rVFo/zfcbc1Y1Rib3IXF3BPcO9cNtFWHgFBr2tErsWPv2SHkJz8XO72EbQmvlVg8UH9Wh
wMojKS9Ywx2NBrVCclBCfGBl+0Sy8M556RGpsK++TjrtlBACDSD+CkoXd18o0E7sW7ntg7NnCe6v
vwci3xw0DUO02P8s5rLj1difz/4dFCG6Kv26npBOGko7Ey5u9iEKrmD1bO5wyEXVc4MJgpZGbWOJ
WFl6iLL2CaBoAK/+UFhvr3aJyzsmNFwznwldXe3V4E3Jr81eMsFb2sTgBhLs/MMWQummyQri3etG
SS9nyHnbjhtDazReyXU9jV6rlc3/IIGyXcqeTpmyqlrKxnxOPFPW0sOQoK0ciOEqEykMNzkhoJmk
14RCS5bCuD6lac4fkuIbyohFTbjR/Z1cL6QLErKYiV9t23Ag2P0KbIsLcijWBDXfPQnEkaY0JKh3
fjxIynnw76QglQ7fXaYfJBWmVOkV2XafKtgCfU9eeH39c9vPz9tRCYnNLCJIGgCGRHZbTcgAdGVN
qH9YeVZrDkxyg77Gqd/FwLnRpft/W01vHJn5v2OFh3+4pgXA4VZXY3GXCaqf5qevzk/ozxByerCP
Dm6oapZNTxhj0h3nQijg3soB5UnjhX9rmKLR8h+1tTzQiEFEeMS9MZqY8Tnty4AYdUBWx6PnbSXa
38zKWtWCoAhsa09ydKuRTFBsyVM0HqDZw7C4vMxbV3Mc9/tQTgSrWQ8/qRi3rfNDnrOuyzh6BcgO
xUJtbE7/+MgZJTscqFA7DDR2qj5YWuRYDRYXJuJmyTvyxxuBA6qI9KilHS8hNrvWTuLdAqen7nzq
S8sM0XOOG9piIahPGSyjY4o258+hbXESP2RqbHRy/TQwspNOo/vT69ggWDXUgDSLCV2T42mGMg+s
/pNIYK3ia8RVDqQZ7uKzHqxYEkY5SwHtYZLVCsF07z2uIl2PpXk+ostNSqJ1CATfoR1ZMZ9+JiM8
4nbgP1YEUuJu4orqEA4EvjjiqAcHIOxTRZolVZymlv6sny+olGUIhPdT3/v1EQq1T9uGNNqni496
MgbWKm1+zJH6DgKl2btofzglVztoyJu52K9kDfsA7HPGlahNTdXxSJuIsmzkU+TDd7/h4P41u4zr
DJ+5/WSfes33XKyhC8QOzVdoTXVbaAmsqw9PpaOBXyjF6R9R7b+l7qYZS4uOi3+apYyhfigBs0fo
8cJPqRmIJOf2FV50eipr13ABAucNB0EWDD4uqzxJ9FgATuZZkkW9sNtAl+WRMmuz+a3ToBozjoHH
H3atsen+nyXdAss3VR/FYoBsJpN5GcpIKYOXS6XWwvkujVhy9Kw/osGt5KlPAxd9acrZi8DlIw/q
XUo8f4GeYedNcKolEpFbJAey40zP9wN2BW0WiuQ8VOLPMy0WskjGbIvT41b5zq+WCNXsF/vQ61KW
+BWbyE625QBFp0yZIpu7fBOmhWIr+q7qUVNs6RGk61wyfa+ZjJ+Y8ZP9tzy9lThdFYzvud1OwU6M
996nVwl39Ayt9UP38Az2tQ52/jLJjAQFPua4TKVecvmnZAtA3eVKmeW09QHdaJ5CtX86cpdXrWMv
7+1RTL+ahszhwAkly0pYgnWZLbZeEPxoldxf4W2OqGmlvFbVz+1Il9H2yT7utt6gpbvthZw+Z8Ee
u9c3GIR+mJpdqmR54QnXyz8YFPRG73t6itaiV0xAhK4NqlFy40a7dGInNnvH1czQElQzGBth7CGR
cPxzClaEhn1Gc6YorSK96ka8MNYYfMscwZCg8i2nSDBnBX7tFdHmx/8ep6+Efh71YU2BzT5p0LkH
1zosiHflllKkE4BemfWFhOQZgQ6KGcgLlOWqrBEgEAIeHkcCSlrhLUv6EceFhfrM/QGsSijZO88P
fAyqdfg/9nPFB/yXTBZ+lqTd83ML/BKye6Yu5d2jIjq8FzsM0BvMmLCLTBgRw0BZucCSKBHuSo34
OCbbRRmFXpmAOOpdKwvptKtrOqcHGCPHDFvVgRFBYsCH27wo8ulRQmlkIttbwj8UmObu/1yWw2WN
g6HgZoOH58DLfrJhAnfUOQhHTwKux7nrzovgYH7Y0eB8ri7GwwHCx45R6j5L+q82fE4+WaYA+Iv/
Oj5XBnDWCEucZtu1AoSlsM0O24bNH8sXEyyJdF8iMHu4DHpYCvDrhMCbsycrhjg9oZCUBDkmepRa
YTEks1QOHTgVZdZK3IRlZsioqd/BS1fKSltFyaEGlSwCQxOuE0n2Y7uDUR1xG/q3fOUXcRS8uDKu
b9tsPnsnSnlrHA2KfQXObZOgWo+MamLXSG0pNIxh/aVAdVgeZ1A3FjYR0J/mEQInLCnVVvSa6Eml
koQYl+fWp3AYayBSkSB6FVgaxE6Gqt6cMxKORFuEXbZzcs6Z7/5PIfOrcJbXLivTK5au7+UorO7z
qIiPQOBb4C9qsrrBCWEEpGdwzzH22edM0B+nV9qRC1gtUTVBU6VY0Sra5QD8ULi6wJhqtBylGrSg
UoIX+Wy/GQX9zuINmbAaLqtqaT/N4OmHqbgJ7pqXgDg0QRMnXiVlHrzzAuvFox7gmFtw/ebFuN0X
abvzKTjwhXs22m3ObsSNekIxQP7UVjAAeJZtBUCTom/OhQo0gieKg4Ai+5hrKOatC47cIs2bxEDV
Sgtwk09lbIK+I7EOLa5jM/iOvCC4t3B67eLV8Pe8/nRJDRMLxNExrb+fNr1oqU+aeYGFGoipM7En
uov1Bva0ioHWFY9i4Uv4YwFVhnDqqUa5Cf4WcN9tM/RMVPwzKaGbysCq44Uq1cT2AdHv83Dcih+O
lLRnL2iiDjzkp0cnWwP6NAVyew+mM1R1C3wHTE1yLWfAiT30EhuzRQh2LRpF4wbPBsv8aWyOh9WA
ioL6zyLj6+JYYZ+N240SZObQJfb/k9BqezK6zajzctekiyMrTKZ9soeA1RnNmWlkj1X/mtae7K2z
eTTN/omvN+r+7xYynaXuJAlKvPrKcRcIbyFWtuaUyt/W2rEm+aWNWn/CLO25S6fAI5jgl8tfQ0f4
hXp7RH4nShXzucSykoo+J1vQkyRcGRust4vBw11DBmMmW1NEKEikvw2wKQwha9ub3szUYXCy57K6
d7UZwn5T3Rfj6kQdiYmpwg1L5mvuxg3z7Ry2UFkBOZDptvQmNpI2qcYaBW/93XEjugorOh8mQZ51
5DJzvZsYdHCtw1yVN17ZKfb89giYHVNgHBqTPzs8TO/aQYaKmjvIxw3TVOzouGBbrHyyGKSn57Ok
+2eAqxnSdjdfhJEieuO7enOu2dDWfuw7K0cLdUhAMClL+32ja9NWL4oqCD6J1m81ZyYObzS0OSMA
yHSWfUnndal3lIzVcjE9+Y9uH2dCwv9QfYgltZCiPQYzy9arzcq3TUWHrGNiFWazRPjvTd24EezA
X0q63M6DAmGvfrE+hEBP3gyJdUuURUMC+tJH/4HOc99cYelIHis+O201Kg3WsUxzpsVmpDvVVG//
X18GmZyQBLbOcTW9IrHabr9KXkVDqsDWQBV/pMTwibSa7v1Ht3K+ir87+zLI3dPp5/RtpBp2xHIL
JQ//hajcWeYOguv4AZdqhV3orYCKF3i6JG/0kiM7wqjHAX9/qaQIi4iuRGfJqR+j/pXWeh8gepZ6
GsrBg53PbD4B7u0khCyZ71DgltfMf1vRyLbPaxsxBAVkDJ6lOj8nJ24BTbcAq17N9kkq5UOowdlW
aACUyGr8BTjpBzrWl/ypoQjhvhHS2oScdXwFloZ2YHG86vLKoARxaJFn0Ra3Zr/2mE0dWVvAd1pM
KxenVvxbWZx1HeaqOeTz7eFYjuEzJCgNsbY3vD3PF6yHlrK21v9lcTQ/honoFdEvelTnOeze4w6V
OCJLjX/XSpp5GlidTJaoqO3mwfctCN5+CGNAuh3gSRUiFftT3yWtfwsGNIyVFDXX1GtR7RPW1JX4
SWEnRA6can9cHHCLM7t4asvjPXOUyAiHV6jZZeMZjupJHej3GFBpF+qhMKe47+xZejjQvVdhmHGY
hzIrflWmvm8Da7YMZ52fsBfRoItaZ3aqv5K4XJhoHN8JBRZt7iE7G3YnVO1sTptK8/231B3WygfY
lL7ueAgcxKcU3R5SkE/a566dSQ1iFSi/BIH2YOS9WjX7xyhAq1mgknYExqHF0+Y9McKBR9G/MUJh
MxEQGLJXg9XmcEOk8OKfxf5dYF+Q/xgxd+46PTX7VZhlvwPP4cbJVEbLmiQYgFdDsap/cPefUrfB
5ZIZAbhp9Xc8zCYUbRh+JGHv9cK1OACRj/baJogOCNuUv3knTP/Pa/gUVuYOTC37jl7LwkyMH77H
k+fxRjNMb9Wkv85iI5g3A+pkjV/Mm+4yTprh6xp28RMLqqlosCjWyo2sHWxxs7+eVaUFUzlHwELq
cVZDnrwYmqmQvBZTC4l+nE8mLjrEJjjbn97gpCaXW7HK4bF6e5oVt9OkMNhvYhs0rwBAbNheIRlu
ZyguWvhteJ1k3hiqnsvWcnf7iVDy+Xcr7aTtPpSAjh4rn78oau01PRXgOe64s+1fNkDbLAzgVtwF
F07P61/xGHJHZvEpo1xSem1cvtnyn5l8hK0qsljonArKWN+dk+swkXafch1CoL7E1HpJpaOFTzGm
azm92ejNbmnc1R7oGN4x3O/+POs2BTayYlXDY+tAp4aS/DDokhKp6s90w9wHYJnT/3cH5ofj260g
3y8YGWaQ+d9ZpZJFwXN6AVS4fS+XGVg0crxCLvdJoBsgifZzCXl6enYkyAGwGToCVHHbGgVsvf42
abZLse7ALPHreFCsUP/zXnBGMtdCt0vxfzubq0DZRg3vjfaxOgLWxomgcuMDFfbyF9KE+4BbgOC9
JsjWRJWv+AJ7DWU2rfstxt3SXQ8VInV7SuUNLeCKjq2lYUnCwWIy5lyTcmxRk4jRy96iIN7UkgKT
l49/U+0/6euiMsY0BHVmRI9vdvZHfob7iy+9BxvrxPV8JnNaypGvj0LPgwm5wYqSAD8p8DpYtaFf
4tr0mQvIbags4vcS6sBmfdcKPXMrNcrs9xxNlepC8FcMkURpOayW5O1CJCzxWoXCmEn2/hrolWmS
kiyKR1yHLBMcZRdGiFMh+7+sdpEX+Zkyz8nqDQyifUgb+jbLTeFnCJf9BTjJvyejiPaZIZkrjgxZ
L9FsgpPyL7F6kravvuRcdnDPZTGGuSOK7YBvmH590/B20qBEHsWZHrEvhaxfqwAk2QFpLTp1zy8Q
qAEw3EaKbDLr7mCAWOf611U91rvrMTjeXThiFzFvzrFBgClYiUw81AmpvZaodqPjusZFCATd+Baz
UoUdfO2YvQoxCB9CTbsHSznlxSXIuJDylfL6nbdhaM8GrpzsoEYGLHwREAbIkP/XNepdFUSA/goy
V6sFuGzJmsM6ECN0f+YVWPcnPsrNYbdwg/vv+i+LXi6PhkQb4+GACjL4JcmpZqe7eOvwi7tdHMEJ
BwmSgIYDeqg7nXYRxFav9dRruXUgJ08xUOezhkL1yEeSaEdDDV9Y0WOEPlHMpximjH1QGGcv6ojC
thx/Qw7w5WmzQj2qxA0MZZWy3ueU4Ck6Ii4r3NQvfKNX91EuqypQR+HZ9Qd6smRaM7iaSCJ7MhQS
EhbYXV2XahhcQyEy0IcLIj2DMd/8ap94bZTB5cItWxCdIMGjisrAd0ZSzpBL/ScPsSVQX6iRloXJ
KGSiK9P82F9jA98yS0PbUR92DVNlzTD9GZXtBSiHO6M4XIuTxXd671r/sUBzMvEOMPX2kEpIV1Lp
38/stoT8ZIoQ7jHkk69Hl8L3+NOFhflNv9dnlEl4OpxHCJXQL5tHPwYy4inzqP0byc8FKtUpb2HR
aQ3hkwzXSGTx6bASCsyWB7DAsTwIZBKhP81Ztz9wmpRD+MQyZnpdiIpnxwiKh1uunaHwq4RN0j2b
ICPnXnMbfabvlO1u7EpD06w61QeqEAlySOoXBdQNjTCg7ucEqk4T1uDO4+oU9RBaOX1HGd2VjYaq
pNR8KtSsR7mKvd6YkGd56Ba1scheG5dTNd8RRVaJUwTo1s6twGZ47g8mQ2KCSUONYRwE/NcE29ls
RHvLBtrDsafrs1St+akBaazSZA2A6R3ZJLdOZX395SBC2SEiwVCAeBRoMzIHSYWvTOxODM52V3eL
+rM1tS7ZB9fVXy4Vk78+aj6XKbxKlpf9txBygtls9klUV1clw5juzMoidsUPMzvdofLUGS/aFQUT
M6sGyijq/hxyiLU8lHb8zYeOdhMNQMpz8LXiGDAqP6WlcHfLPVm3fVR0KhrH3OszYcpKHUbV+NwP
jxDGrr6CBP8BD1S2yjQUGY4sP53b9IsauVwodEy0jcg/tFyI982zZgh5guIf6pWHYg6Mz0Lm4THD
EbWcCJ3ZW6xbNydUBxWR4PO4SleZtzv+EzttRaCoUOPgn4BWtB9Fa5U/tlFB1BWMBb3ZhHq42Iu0
YLsUwl9Wq3L/L1NTS+kber4AWl5yCZjK5p3xnKSUwdVnQ145zxxWudZ0qZMQhkkm2KeAIeKtH1sr
TGwAJI26/u7qxSI5QT3r4H2OeX3ilqqFfPyK8y2SG7jpZv79zvFaOvAXzubiIv2rYPfwLV5J0ORl
ZUGWyB15vqRA9Ha2Tg+hFTHdWwwlul1Y/22A49eZ8/y5L0FITD+DPAOMdKzJ+rQXnwu+vj+h29LK
d+PDI4JzkKComnCRFOFOxdi91mf0JbkJbKZP+8MyftmxSOM1u5CfHutGIQ2xmPsE1CZv0duIpeAO
QEwInsFrfvicN8Zc6XXNWEcV2LNyeFXVum3zYzA8aPRRESNz4XtlkGER1NZimwo36fC0mjI9vhPZ
xIVHtL1tgumt/UA8Hn+GQnZtlKJez//hE/CALTk28pBTG3WBr3slsIkqlmcY1M1v7F0gNwqS57yI
FgopFa8Nt1qFszBkC3oO3Bu34xCem/B9i3djJL3OAaZB1YLj1sHg6ORR55/rZyOqHTfeat+emPs9
mG7a74ErrpatUCYWxyCrhloQCxnR3AWY23e9d1fq4zW/+Ox8KKoVLLrEkN/SKN8zrj8a+98VoUFd
aTycE00jYV9dOCzQCyQUdQX5HTPea4KTp8KGTEqUXptoYidCKwk098aMWzdyEVJf5NCBmeh7ax9T
p4yzQE5W3cNy33bnRreN2g++TLyW6E9Pt8C88MVFwKr3VbWZ9GTAsZL/pn2bc74Vjal5JAazYVoe
QgRsx4q9oo0Yi50K0AwwAfTRjBShIIiPjqRWt/cGzN6T3CPmr/LXWWP9bBxqAdHp6fbgkBv7QqEo
dopLSWNa+Oc85r/BcoDFEJ9ei5RdeRK+OWqm6fL/GBY1CSPAcWdHB/zjFBbwRiKWnivW+DMlSwyl
+LZS8J+DK/K/bxn3WV0yirL7yfGy/cY31t9vtfExjvRUDsy34bsWwLLMcEDDrowhn7O/1zJbez7K
Qr8xt/Gkb2BjXwDw2peJtOMNb97VAdNMXT9Zao91W7ECqal7TUZhMkb+fVFXGmcrW+La9dfF3KhC
UNKkFBhTCtsJOvKXOhedi0h0hmsRRYHhvJDSNDMQFwkfvO6bBpsRi2dMHu9sQ8WzwSMG90I6Tn2m
UBG9nQf+AaP6yVHz3wy68UE5p7gvEks8cbCvVlJlxQsCHyEwHxUwqoQpoQgwEnbFMJZg9JJBZK9i
DX6eOdLZpEc9RVvsbpmPPS5xPVsWJyk2mCKKc5O1YcTTYCK4bHrMjbTzoyFKRgl0XPtOY3uNBv6/
f4Iuv3wzVWwKdmK7FjWQbwkrG+gn+ET0mBdPcR07ZYMcVN2zOORC5RziLxr1rbdHd/3HQjuPn+JK
xTKiX8raOXNUsvvBH2DDyDAs56U8FZELi7joFuhO/ufIhiMgKsHFcQjN2mMVVxNXtISRSUvscvRf
tssy8tJs2Ep3Yj9DKZaMe0QQKVC6fTWA93CMwJB9/AJJFalloWqJ1DYaHpMzPEafoptbASxO2HHs
2ih2qxqJz4ClBdeAB57eqUFvxDzhNgFB5Y8c6L81euLjQ/6ZEQoegN+kpyXrx9dnnTVRxcKEXu7M
v07YNwVefHh3C3BUrHxBepMGrB9dGUwXlRynSAnTanwEJLhlr8N2xY34jqTIsNiPoF6iosJPqm9e
kOxHTusWDYnVit5ugtvuLqBwN3E+bMV0pFBv0sc/GS86Y79RQd202XSqB+hyxsNoqoGUFKGwy+Kf
FeCiF+x/PFvdQiOjWGYN4ixHUWl64VbvYQTm4X6VkVDbJx5kvNYYE2r12RD9fmy/n2T+LQVjBnpq
OGptQtCQD7lAWpSJtDeHNi2z7voacr9GzvcvnBaAtjS71HrZqzNdsKsWAZcOdrSgo3BVKcQTM/lE
VO2Vk4s5tLDJDtix6KElzJz0rg7fPpBi500JWPolWScVll5xhew2sg80Z+CE1dlBFJ6CnnbJl44q
FCczn7pKpmhL4euB8qJMZxWOVzAedpQgAHcbSPxroTzZrUc8UPYnQofpH7F3t8bvO6JVsTDlaon2
ThbgmYKptgIDKkO2sANxD75tOV6y7h2xl/Bq6pm6a8SZtKeWOcwQuCQ0+7dpVfJ0n+BOhfLDg1fh
IBQEcXfHqOSVM+lv5ap/CrXJy76Qrcwy2kWy79e/86piKKCETf4cwpl2OLPwanBKiOouX5t6KUrC
nOcwBe/18J7J/um2pkZ0vTB+yvZDnsHnmu2/UMYXIH/iWLtTFsGHwp5ZqjT5UF6frVURdbuGgd4n
tYuHvypTzG8hnjOQMFzjppANo5ikMRQ7yFgtUmHQxfYSMtCPUNC7mZHV8oif3PkTXQYKIT16ZJV1
PIbPnk1b+UOFbx4PmdlsytQeCHldrl9SDcnp8adgTnXFfc1pP5PJ//ADnoiZ5GTTAg2O3R+NwB/I
kiSpwzo76cgasW9rrBxz1Qiu/+wcH+TUQlEfIgUP3jVUfdc0+mi3Zk+waNh/R50EhN6u2swSoYYz
1CjP9oRIvVs1VTnLJwqu0mci3dkWhae6+ifYEvRxN8pFiM6wBpKOFV4duAENKe3pI0CiOx4m6ccZ
OTqMP6jteZ6IEupz4MetuhKR3wC2LusaGezHK2KqEEjUy22mun3oL2Q/sHtf+6UGUQqIepiPu+Um
ssmxRfRHllSw+uCN2sfdaD40KNrDO5OI6tvOvSoPdWgc2KGv4sK8eYOPBzmKbY5Af/fEvYiBTr4d
J+8xrn0muGZ9zHZu8ntu7zecqs0uhycEa3QrR/PyPuC0qS5GoVzI8wueWTGJq3smC/gqkKaAoF1s
j32mld9SJgXzxrojfTUqke/jc6uTY5qWyPAPwz5s9X2Y0guOg+138oXzd2+ovTJktQ7F+UpkKyiT
ZB2jTJh72t0cMBgQFRg0G3tqTyPa+Kmyc5bnJF6ARr/LHOr/cOAxydDpqEJcPrzdlzSPYqbgSb3k
srY16Da96BwnXoHbY5iKtsYqQjEc5XFL7s+BLA06uIyP7JG6ymJx0uD0V1Rc7l6W6YpRPxxc1Xbg
gm3FQJ2UgvnBUWEzS9RF2sqp/dJGSiOrD+JLX15gBiqDXTWpBHKl54Wdc+ENMsiuHr/6434IUJn3
IlfCya0GYryupxwS5eMIC83rX7EQC0QGoyKik0vaUOAMjxKbCTajiNzryPfNg4dAM95l0M9/GNnH
HX46nBB9HjpjyjTlOuPr/+u/gS1s0n7YV3cQ872LFp4J5KH7NYTzYfLmsckOVnD38WxKjErb9g6m
CJxTMmD9J+r4ixhDxY6ZXQ64B8d1BVM6JaXHW0fUzBmXN2qk5XxG7cCCUzbTuOFQNh7KkuHsdN9T
UMq33rK9/kC9AtnmXwFMHMGrn4+iMuAh/rpPKT/yHu12wu3fg3x4b13NNPs0eKkJ18NSuoQVfk63
cDu98burrRmGA/T6N/kpja15Ak5PdFOqXH5aAbcK3ywNbSalF/9Nw9PMP+0F5GQ2LtU4rtmvaHtM
PtfoYlXwSNRNgqstpOobxp7i5bU73RwlPDzZds3vYACQp3m3+hKPuXtE9d/F2rFrvkFE70+6xiR+
5o0SpRw2Ww2Yg9Qr+v9tOscJSFbIWhiDQK5zWuoHzRc7OkKOadue1rIt/Wa0vzFxF+IX8Za5Gu9N
wStSchAnMSqbPN3MET8uGHEB5unqvKMGHNvqsZHHdfFXQUeyTkZ/GCdrorNM9ph4egKKpKD/LFzJ
3QVHInMYM4Piwe4l5Xy5j7gAe28K0RxxBBLiSBHFju1lQYRkEyCiXgcGGn4OyGtRp83wwxH4mxtq
fbuFtEZ80dGAftzb/sfDCAT2XcvKuphMTn2ZFkJ8Q+Vw5GJJJcuThsMWkDNyO4keJepa5HYDQoMM
3m10RiSwayezCPLUlsTD676jcOJHW9QoBUJrvkDuzY128DTG64plLzpy0UXuo9r8f1W0WmZNqpwB
mBOqVJqLO6DXoe2MhnpTdm53le+RcbZ+grS9PDYmQZCdiO8XMDnoXkxD114UCk7se/3PbRgf+PCz
RMkvFYqwnjlckel+TkWjofoKuomwn5s1UPRC+fGA7YpfDfYa/FaOMW40M9U7s+FZk9uobwjhEsg1
djLqzrQFn0vSJjFpQaKd0257yJFFRcR3hSyfzZG4TN4nkOxIBovU2tuVuvZNkR9hTRiEEmMlY8S0
bppIhZZfDhYOfk5OvqMmyuUnt2n0X+T38ZuIk1d759G2GMl6I5EcVXsM5+7YxCyssvUooNanJPBn
+SLSpopX4tZ0Xxgz8djqqAer1xauUAmgNxO2gheNhe0sBq3JyughXc2bisi1uyow1pWW6zm6YBuY
y+Li9ahK2tNUAlLi3LgaYjnywoO+vFdtoQesJMsbuYwlyj6EeRcWS/nRVH4ZgbegB9e1aPNe0bGH
QFiTyQIftz0o/gMuJ0Gm9A+COtBI3PeEMGzypsc/Q5mZH+oyoq7R49YxwkuwLGaFXgvL/fk0hvzL
Jz6VFQPw6Z63f6wZsZFmj08ifv6s1P+pI/BgCgU2hiilWbHhMfWPgPWLjfY4PfTI1HJrf4V/NzbN
5kr9xlUzUrFYtu7Ftc98zLVng6eeaF9iiZx8eO5mQ/uUSvxLSWsNJM1gAI9MzfbIkdYSDAbSqFUV
edu/S8JlbR30j8HlguCPaXySlsh65fOiwEtWZ1AEPtJtRqTQ5/26eMqHVdFZmeF0lm4epjxxlblu
pC+nR082t03Q0uWecOsXN6DLJM82cn7q0kJt7GPRqz775RwAKfVENOSdTjOl7io0DXT8G6yWmb8P
K/sD06nzfCuEvFs0TOm+ZF6Mi8uaMWcFPuDFvSXjoTpynf/kDgCNzSnzB/VvD5tUpagjrt5+P8h0
nJTfY/cWMAipTnz9w9pMoMwvugwcajg6VbZsGKlQZy1KlTpe8mu4rZHBA/FH4IK/FYTzwJKPMKl/
iCrZz//m++I4HZ9VKiUac4V2pAXBnriS+HL8UNvog4LrNJCIdiZ5Ersj+4Y4JfQmv9CfGDX8R2yP
eFK1vkZrlmiKkfFjbuwYT/capsN2mLRYXSNI4zmg/kHYhtDOxfN2fTimd8a9CtVvDtl18NXYlhvJ
S7/ezPQ+DZJapGl7r92cJSU9ohTuuCQS6MsvNFiJ09XT363vSauypJiXipydv5WmfRAhW7jEzQsM
kq+Szu5CL3w1q1iDs60BF0rOBtWbmy+YIVEWIUTTz3gAXOIwti/WnUUDrhumZVrqSuq0cAi4bGBd
OuLNHHEgXf29Mtg/tVMSS/HpX2NRUF0YzhkeimMMRm3efY8hX/bl1ZtHwNhRjy8+eo+tu1wawDpw
LL/j3l3DpeMPfAosjFnxquQz+/WGXb/rs5r2lTm8bG6842QYfKerWLfQam95ANREqhbr46FEAcpu
+rwMCVC0K6NWVwvAS2wIys7pyaQRs/bNbU7+V6zXGd0h93klNeWffxDFhmjtCeh5NhLGSkv53r3n
gDl90k9XhiDqwOJBQ6ckptQTA2hcXY0HWM5ggEtU8Tu2wedGZRwMVyXJGg8+kCYdZPSR5Jqp7CBt
g1haaq/OZfX9mTKw1f3QyXBN6ExPhCx02ixNdWvXv4Jl7ceaOIU7kfMYWHb+0U4Iopg6FefPpAxx
Z0JjOSJx9GFkCh8tkCd7Ij3sr9e7eZVwHUGnDz6perZrQqrwr8flEcxr6n8jfunAvsn3/dCOWRnz
VHI3er5pHWPi45aZ6GJd2OhOjdBKnf06wXgPi8qk9InWAKWRDwE7Eh6oLJmV9txUNYAqOJvGT3zg
K2P0DVYsPJlRYL7VXL3ObxMKHIeKKG8zZv5N5ze0jJaFL9A2QHUzr9G27ZKukMmSudllBgkG5bTq
PwMeKaLm7Zi7bMymakhVC9O4AP9treaBzAjIPEPxnn44hn0aPntn8iakdcrQo2k/DnBd/zaXI0LW
DJ0gB8abtJHA5084zhapRFWd0kKCm90j5OKx0QZBrLiZ4JeeSn3T4QYkikUaH0iBgSrENycTILeV
WEGsw8kU4CtgjImC0T+ooivAOXTOgaHesq0lNvnW5l9qK1i0xOWux9hEo92mMYt0VFkeN3/kr8fY
PP5IjNA5Pwb0pTfL9BWPsBfvTA+0l2bG0Rol8SmA5+LUGO06pf1lESv32Yw9Ma0PRl4YI/FLdWxN
XIDNshKOa6uhshZJA4FSwXpQtn28JjYkZ880YBkpnLXpt8rLf2ZdAe9T5UV3J+sVaozl+4HTPLtH
uKoKzG/0QugFHwwqfRkcxybeQyxnpXYqeTjB/Rt43aqqWncLP1Z5RoqY+PSaX+Lhr2/J3Vt+3i1W
wuQByI10hQF9H2/mGJzgdNuScLiK1HoSSYT6ONL1rpi5HQTBUo53mJvJTf2eafQgooDrAn0GP2i3
DMWQJxolNDLYnBYrqX2pM4RGbI086U8r6dsnRE2agFWzseBbSpGXrCrjpyzAvl/3h+6CWDQNVJ1O
gAyzLOApXykBwPqcYu9a/zl5oWk/i/w6Thm4nN0M1mjMK8xkBLEkP6YjmkrqZhpcJ+aPVUb3V+k7
t02S7330B/9O07Hu3n1ZIJ1ynDi062WwxgF/zP70qytVR58L/LR1cuHm1Qt6zX2hiO+fJZuP76hx
dKyEoEl7Zdki/5dLw20FgZzM6carL3yDjf22oc7o0+ou1goKlEjt968DCVEiC/M+t0I9WUDS/4Ni
SjAl4Riz6Yu3qN1r31jDC0+0JgoP/wAjMly948xulJ8CPe00j+EjLqGS8XI9Rrpqbo3w1T2Qnus5
jObhIYrNOWI/z0npS6t5DptsoaAwITRm2XKkfuEyYuxNUQwY9SRLV2DboLJvcfG56Td+c/ZeHupK
eKz5agGWptcJDEMN129s3x/j+vsTdeBcrqy/puzpYWAEfzhm86VvPzvT9a/UjjSCAjgW39urb/RK
t4qq2k3j86SM4b8px6zNQcw16+cjMTZs2L8tZfwA1Fs/SeGYhD8rxO0VSfcsF6bZiYjH8s8KET8x
tIWyA0UcbxJ7sG6taoTAgME6bNJAItW3470hxt+c+HSef6e8gtujVPUhxotKkIxp+FdQ5SUEuK/R
hAQSupKBQwkBzzmLUO1p5zJjv3yF7U04OICHMaX6hJA4/wKjeKravNTn2U4WAzFE3cXgFYQcyzDL
0p4Q66ynvaF40YjWljUHeXCnX6n3O+w4lpTMLzQ36pN+tAyI8HIDNZP8z/tufbFw2Fd6I54PFtq8
bm+2QuhpaYblyK5WSiURdnmQ+P1L5Ndc0YT5WqQvHVUVjF0WkaRz1wpcAh+pruAiR1Jzf68++2/N
/vN5eCetap3D65tk8JCBvA+FvvFSjY4fmPb03sr7RaPcNxHXohFk2XNU4zkq5S5HiPGHQtGKRNkh
nOfcG1zipVWBNCGU7cywwEdHciNUh4Se4FOqMBJz/Sg7T8gy3GZmDs4EDK5Vnyku0hQ4DB2z6q4u
t2jbGVOfWcLMam+k2LowD5MtUC0M8rmgfFsx1NnegtWiU8L3UGXuqJe/jiOnVRI/5aqDj4BwSvzL
FABdGUuRL/WcDwLDdgImWHvEQ4c4ajELOenGqKGO/rUXGs/B/SJmMwXxcgUALZhoLHCcU42nJvR0
1X78/nVI1i7AdN1GoeLuyewBustxkYg/txj5zHGQs//fWqm+kLC3/YCtS8Q7DmxT8q9Wq+QjBdGq
Sr+Y6+Hiy2b25gWxu6FBLk67M3v8J8s39UZMlN29T9mAgn/QOK73bq5BlH89Rtbmv2R1qPknVfEt
jDvM/zxZbs9+c73cBiQZ3FaUP0Brxgmv7hHNYOcyNTxwxOh4Ag0jU/G1aju4kPpWByYuBnhWZmb+
EWGYVvwgD1bEajgB48cz/2nAyDELBZX6bRTg8T4ws/i8nUqJTvsKcWyeZRwEIvoecHiOJo7H3zgK
7vssUhErCELSEoR0wilWoB0OwN14MGXLM7+3u9egH5ROGvLuygMh+bENj9mzRsDC7pfEtRdbm+mJ
xKmm+hLHGSD7iyXh2KhQTxznQB/TCGfQUKTvp4gw6uzqyoDq7QCCb0IzYf30EZ/eSXY9A7/85Ico
mB3p3CaCaH2TV5vZM7qH/0foJ5lGrpnADQKRo44CsuiKLIcb3swJoPg4ALcWQnCHW4IU2TJcUUyp
ppmyDWKaBJnO9Be8D2gUmsSx/2QgUDQZgm3p0fXLAkLVRb+E0HfJs2eL/QT6NJv59IpmteRYzgOw
6m/6qNZhFCExDeqymjKaAZ2/weA4BYAii79rZCrzZANjcVks5rKuQ5FCfiCVN9ZTIer/aB3gjn7o
T7xTaOUpGj62pNqRmK8yln2JVAWuA+J5q8EAxOSB+oi5PPXpVhDshtwtm00hX35BuM2eUfxRRM9o
h9nOjzekqVVfa+1QKp0+7Qc/g7f1L4nxHTchMEs5PWX2VN4510cLt2hoSk4kCIL/KrdeaQEWzKPY
Idwb4ogUkELMBSNtp9Yld02WcGsWZvthFK3bwoY47cQprfchGk/RhC4EGkCj+kzhcieg+3nUn+Zx
HnerLKGdudvCqNNg2mRNECEWf3BR2NmQO1gmzYlaZcmyDFq7toZ3nTzuSK5vXAKrJQFvBl4D/xDf
/P9rJvCgVfh/deX7WuF8/okY5FxmjUSfX3PzxRS3d4U8BQaly07YqrYe22qkOOAQhVRYdiheANHr
x1MlSnudbZTO7zw0Q2dYhTH8zM89UDrUv5poX2p+nGZlcqy2EQ4HJXp2GgmnJTtyM1cA9XOzga4D
fSHRUtgOJFiHTJb8li+4eyYSKmmszB30YyqbmRAZKTtn83zvQ5vJDSnoveWdXmecr7MGO9oBBMSh
+y20cSZYVNKwhypBp/YTAWKNY752ksTAtoOlvij7EUQ8GmsMLqp4ms+i+6JcYCOgD7Llupg/ks5I
rWFGEsyJKqWAil0fqIAPlIW6Dl3seSNxLzu7fmntVCThmWt3UpPCmpenC3i57dxS4s8c/qVOr5mq
F1DxVCbycuSJ1gXYjuVNQOPV0cz+7Vp89z4RoqF6tBpja+Vl0yvE4PJGvOfD0HaCtxTrSBnW8mpJ
s9f9sbR9X+YPjQxX1bpHlm0WDbMPuvtiqQxaRuf7EqswCQp7eB9wUvVH/oQtvOdClyB3YVeZoU7F
6XgcmXljTSpisrwhn+qlNhQrcTZutAKnBpjdg1UY9zrSbYydL65Ndgn2acKVXCkyIB5zQGToFQLq
AOguvGbIiURguCdPWNP+LCzO3ZCM3ZnWx8p0bA5LxX22TzCqHQE800fQihfT2yB0jxVBirSjH0Cp
WvrO+gbwa0Ww0plwYzCNdOZzrm85sacr9dPabniXQKe8ao51oEZD6eRpzF9rfyHXw4/IXualbPJO
tkU3YAqv2Oc466yp4llEWdfhI3vcI51RtZJ5sqCCXVp1u6RIYUcjpeH7IXfwV7OxejXC6qgXV80b
aIh2Ubzbl1HIx9I1Yp2t+U/WY9zbftMZqpaoUmJfPyAa9V0JdLQ635BjvYg1m9/0AvvmYwI5p0tY
2iDLvcyRQv7Tl4U6A9KkGMf/UKhhq2lLvUT18tm5xOemxHBoAx66bYYg40EozNv8becyOKoX32hJ
A5cZ13Wn1cfFLeiY3aUzQv/FEelC2BdExapZnujCwFHBPWugtqKT3ZZ9TzbqWGddCUDaDFVbpU+v
3t7xOmRh1WJalpi18oCIApZu0nXLnRS/95A7kBlW2kWM5S77HYYe0Vr8nxwxjl/lmeneu7bLbf2C
Pxk2kZ2et0Vzdvo55EvANgTTIHpEK0xyRzKoHzVpzNvsRhje3QoJ7+CTGrK3eeh2Oe+S7FBYYhhG
ZmoMiL+CxTDaBRauq8QamMck+v+TcS7t3NhBlpEZXXeDyadgQ75dPlzMdt1WtQpvgHKnvb1b9FRZ
X5VkD3v1jHjjTOgwrfWWFWKucWIdZWk4WD2bBgRffocXc9gOSjhATmfNkkWnryt97ANgxkzfYO/r
6+CJpTpCg89mjrBcYSdeze6502TJ5bFjsj9s2/oPmrHuCTf6yRYFXqhSyte2NsCtB0kIwDd/k9Vz
iwFWckkWi+9kRDkfjGIXem0mFgc0FUc14I9PjsE/+1xELuB5mMxipZ0Mre3qNLvZlXS1fXbxNHVa
XKkSvBwIT5OpHDlhbVJW76+fnwJCA70raL4s05RZLshBZ+hfnxafty1fADiHoIN6cetZWceHkB7b
5ec0xm1vstkO5WeOgbhz6UjWTevKHq47ADo5F6P7oW84JkLIBSwaScg2EcoWgY3Eo4CiHwHPDE57
0OR6WPe4h3jnh4bzQB5S1iJTwavws9r06vND/0H2wb/03oKKA+YHdbxmEQzoojQUdSx78ijr6LGk
iRj83CPUwr5q6+vRyGcc1bHxcHG8FfaxLmrU3mwlqQ9Cgvmxk+JkC06oiV63wf9G6qQtv32xd2j2
3BBF3LqEgQei7Jx/ODLTfvLIIizPYL7LoNBJalGTrjEWLkiGBIDPOO1JediMJAaKPHAQuelCF33z
QGHK4VwouRTMbCUDeTq+Xq032urJ8rDdtc7I7FCYj/ZBpSHs30eh15aYWx86vZEhOF677771kLtN
baCBYJeBc4+cSugi/ivfdV4EZu7az4a2NvEhqFh/MaiV3dLLt5hdi1c21q9SgFpDL8bO5Gh2NJYs
/seIgdNKnH10mmXxVLla0amWrHlIjbvMQWxW6ld7sGgyhSDg0S3be3F/o2mwpTDXrXFmjNCWjJiE
7Z/CBTkIHDjalmQHrckQkRH0/N0iMnq8CGCkFpFiUfOjOzERWwSVbhHG/3eWARJ1vbFWwjtqq0Jl
NuslKmB5vL/tv282b+KgKJNJjwm5k4QFxiKQEgASMUGOLoJnfUquoAJufpPhZ8Wcw/mwZAW5RU8Z
+NzZdQxZe4ZqPHlr6BtJoqqRRgiSWHpSydCwTEMaGnIFLN3GbflH6ETgyvupe0gFEH7K2qY24fKI
/vxm2K0GvImLIoaO4KOQQcLGS+66YyObOWewvFmolwiSfM3FB7MzLBtQT6cCPFrEbzrEjq+W4Ubj
5ew3EBQj44ZSCwtkoO7jHkSHS23VkHblGpfs5oYD5vTCay8S+YDgnwh5B2mYRbWMSR4CQUJ1uy3r
IPEs+DusOOJyY49TvO1PgqMshD671IyYP9g1J2F2EVGttjz4CktEIo2TKOUlQN2JzfCHShB1kdUw
acJBXZ3cOY4C9k3v/6RzIOtx9b5rvUJQHIlrv9YbXUUOjk0mgP8tMhOsq8xCsBXs+BjWBFOeg3c4
W1qfGo5MqK2VawSAXZr1XkkhY72rF/Tr12kxjx+/Zh3eZVQLruirdP2XABdGpS1mba7veFTQYK56
D6wOzYcMSfZ4EO+G/a1oYs5aaSDs2xFO2ojDBhUY6I1VVa1XNuOBi21dAPW/+el0Mzt5oo8FuurS
o9aOJu0qdBWqu0femZ6msdL3eCgSX6coZX87C/wuugi56PsZmbc83udBuYRVTWyhsJuo9WVwzZJX
qPmnG2C8664ElqHWnBA54LIKXxmpPvzxZHOeX1MrSBRuCjTxSDb7eaeFdFJOpWHw4sN2FS92/C44
m43fzQ8+9c4MeY40A2GXKH2OgJahrkduBOXynzgPp4JzsSv4O6xU/QMRp/89A6NtmP6UNfe6DleL
35cCnppUQ6GYFZ5MLH/Mch/6pC1yrn+z7Jb657cYMrNfrP6TgU8E2gtWZt7vBWVT9k6MkjRNWMq7
hiiUbFK3XA2a/d4jrPffldfToQyzhHO0CnEpILY3TmbQRC8rV3vTryzMIk8etGvWsykJ7COQyP5B
6Wo5ld5NeCOL8Jd372KL5iXwZe7eHtFk+8FhAjpvp+ercrhohWyK5vcZ8QtOk/lb1vWOXVifM77o
MRMjFwylwBsDCssxhi9p04bX1HSEE/Y1h9S9qpClzCIDuXvPJjZ02lqKHlcohPQexsBxKjnBXOs3
jhbCnnlSx1yT4TosA0h5c54pg6Cx5KQiHnGnp+XpTpR3X2wI88VpCdMrGR57qha+AC8jWGiBhiKs
2v92hdE46NE6SLc5c/ltSUAHvhgp1Z2Q3jgP5+aKoWlom6U/qY0jkPgelpyRr8q+rlFq2ukaTRX2
WMn2HMtkSTDaRFl+XHSRhXJpU9hU2t3QkxuPhWgDTbXvE4khcdrfHI+U8KmMw1XXf1Xkgnony7qn
OlnwzWidKY8czFW+cp84pjvVTWTRELWkREOwCbB5CEAPpLwcBlxzYyTo8bi7uwof1k9LznFZ8QSE
6vE4bXf7zYPCZ1/jWIlrfBzSfcJAPw2fFVbUI6peRcV93XZE4us5Oi4Voj/Sv5x4nX6FJMvjJkDg
6w3ruEY8JAnt4T1HAR2MpgJpU2k1QEjorc03aj7oVxu6nCJWV1lnkB/VkZ9E62kro7jwjZXtbbOd
uVojmWTLHgDLkztS/K43V4f/8DGCBVMDNH3PWkjbxTy9NSRLlD+CTxtu8bMRdZtw5eQAQCdXCYpc
55bQr4dWq7hhsbLa7GO1r61/m0isYuvdJvexDArt2NCVdX5uQP3ws5XwLTnSP6tHAE1m8WidcLkQ
TpbSCg2j5vUl9u0oErlm98plu53w7OrZPwn3eovW2DiT8xpRgYfAg7xGJT3t0f5NYkb31oZE9Mf6
RBImlAtHgmkbgHQwnF7r8GDShIJmV5ysHRbHhuP+2e8IkmbUfQIoBRSZ5i79qzex/2s7Dp0svVQh
JzC+6oTHCgy8sIiFdxTaZDMCMEwAZYMLWT3VmpCux6waAI4A4P5gWcpQVuaDE4FuxQL0zaTk7DAV
U9fBYRXMkBRBkwfGhVZbYc0kD/+xf7EnvkIh0WKonLlDRjNYePqTcoCYFmcusA+mU8OF2eR0kEx0
BI+ocWbCEo2GqH2RylolGB9ucfo3mkTed0qqK/EU2myKRMml1O8IoB5Lp5K9Y5D7VMsFbHqqft2H
9NTn12R/4HZF1KTJjHqt7gKb2Px0niNYY94rjrduvKeRNinojerM5ktgFidTUyabzkLlxfBUOUn5
dRhnfgTe4TrrBAd+w9bF8qvh+HTrcxp6BEAwBTwhWrkEUQNf3FqS3OzY4yAEpVBzBc6tHdFDN1/e
VCt3kT2+rXQJwSKEpO/FsORG5gl10EGcTWmgcBfoGe2iysCKo+7Mfnjv7jd/MWgTXNShSEiJKaHF
B1fqCF0tfn1C0aU13oPXlW7tFmOzndebGu28ZthvrdrIfOCR0sbHpJw77R2/v8ac/03NhcbkJ1Q4
PvLnSVsK1BK6u9IHNMBL6Ohgonkd/P5YUYlr8OUVQgwLM2ajCNXKMx7RU68QUCYIgLCHTvkCD8p+
z54GIUnUF/Pyf/6id8qCvn/AwE/9KIbM2/tW5mlz5O7qEQNmhSn4fiLXtH4vEBNRp67WJx1+E4kC
1G17eQ2p1I2A1IF1y3kch38TQ7jAPwbcSHNITn64roIBA3Pa0roQ0y8+NTTa7YyhsWZw25MVZcER
b0Na7jZBXuP2MFeuLtEtC990CB3JkR6CfMelvOiOry7U5M/pzg/g0H9zXPQDiyHtjEU1dvUCI5+R
XiM2QirOh9sGe6HX02oMukgBumSE3u28rI+0m1W2TWVo/WbZ+guLNB6Ux9wVC8AkMZ1S3xBdARDY
YA87XrMxEWVEuM/1yh+WZm8OquloJzvDtAK5gmkbAJNrOeqABGfTMJRmZLZFEYrXWyh+Of9pEtxd
fVQHjxSFtiDZ810TtzZ42jDwGljs/LZEGQ1VQsKzkGe7apS9/MQ7AbtuncsOFY6Us31RANEzWpnR
2it4TfLBfS1+ppHVNW22sU8Vm8L38d1RL6GFwNmbXn5YZC5UGw5YsPmLq50LZ2H/4TnUDVQKVy+x
mMTy6ApWjBXJ6sFTm90yHF3nMlHkqCkk/hinys4/fVwKBtBJD/sGPKDNnuPXycA/bpqRIkZGniMi
PUHttfep33r6XCrcm76ZgTT75OWBe7oxeVtAv4wHpDmy7CIWnk2z2gJ374IF3QBBW/JSXjiUp7FS
tvQNQUzPnvBcULovhu2wLxpVIF1pYOI1ne16HYPJXF+Rlh8pfamUV7SXH6OR73/hzJP8XHC7ayTC
PWdeep9Vg9dBynMTwfltvBjXk9saOwijoDnQWlOmHFD99eO3DRDJRhQl5r5IpbX9Aw1hZrdq1TfQ
8el2MS16pHtSBtp2wAHG0Y/ErEhkdwO5Zzt8kMQsWToJCts0nB3PIWbtAfEN54v2+BgU55vsUQvT
clr0+We+AegkMirroEZPtQc3kU1c6p9Y5nUNKJ6b58YrRHRMCJZaa1bkIX/5LrK0TnL4hnEhWTDm
uN5BU2CIMZMByj1GsLceB6oe54nbmshTadIszHiZzWcZEc+UaqOybiRhbVAR3Utd5kYCn0QpMX0c
/K/06KuTpe2baydptbfVrsxu8FF/Sqka2eH7aaJV9DJ7LANcFAMougcBHGKTvL2h38OCh29NxOmA
PNR+6BWChSPN+5GKBofVYhyiDrqHuR+Qr1hhM31o/Hf+cIQ3zO8YhTKjhGlRk/fqxQEVTp/mARSh
mc9INkpDrAIqAW56YVEQlG/EacyY+hQvVx/qkspWyZHaAAdFPJmfOW6sDhe/tCrpskSKZ2FvW2sc
k2mCIc7+SlJRPF3fVjmDEFwvHv2bW/IGbAxLCxwGjpt0q9a9x3epUsWqU9V8dUJ4/WxCw5MsAwCm
RjTqtELjSsCX2R3h+mn39yYDh9RhOZSqe+00PUU4F5EFW891J/ZPBZnPAiHIfWBXEKAZIsFZ07cY
IjydypT3UU6Q0a1d3xS84gga/Gx5wnsZh+nsGK/DCk2ybZuWzPX6Xtl2u3XjVGlz4YQtPhgy9O59
4yhpN53Lr7n0zscJ//aXI/aZ9zPhb0mm2/KLlkvYYlQKABwhmvnDBoNmZ3wyhjF78nTAqWH1eLFC
n1rSdJSmbk1b9gVaPLdFpZ5V9Tkdr+ZR4j/78Yi1LkOkjt6Bd69xOXbiWxdNjffkTUBTXo8/C2oE
/jL0cK5TP3dxCtjLN7hBjr1wUfNhf6UeD9RBr4WBAGoTqdgcEe7LtHahWB3dXxqmBRi35qzzqQpr
cChT8y1vqGFlKBcf+lp8+fzLSLOjNbrKCDqooiMNLLLDB8YBrismh9tiOKtszANBuqCFlVewYd8g
7KWbC24ch41hpkaSjbHVvnowWbLG7sWDnBQSi7vpyZrf9xKEzj4X1bhS3y3uGP0XUEaSkM+X41TQ
g6EORc+WTPmkhaAF2Ne8lpFlQQwqYGwouCu6Ry+D9RnBr6NQD5/MWhXbt7wJz20m0WCK9gWpPvKp
VYxfZIXWuDEw38XtEubz/VclQci9q/QaLn1lBfyOb/9Rg5OKT/MxtspAQT3/NAP062IUXfDnOxG9
V5jaFo7tbHlGRi7mJxI/0JNc1034p/gUkl033yF/Oh6vF112Cy6xFAR8mUtaO86h4eAjjnCCAuXG
mGkTM7Q1ZQhiR/27QnII5Pt82aCRA0TgezHMHVV28v0mW4J6eE6RndPusi531pQXgIGklQjUQzVi
Rd/TqYC8SnoBvJ/6XT9zcOygRPGO+IjvMcdhQ9+eFUlMklop9tg71bpmengz+hCBQNi16aMxVG06
+1dHqcgciPdODsadD2G7XYtCp37aJBIJF8Ka4G7TsHLUU6PQkaiwFZprTUAPGSpAArIwAePONelR
Ls/7lpl2Peqn/hGVU+mg/5sukbKLkx/XFR3CktPp91zczAV1/3WsCbVCFm8bBXK2q0ynggujrbHv
Tc6vGk1Qc2qmqq4mLssh4i4JkazPktl8HQ0ncX58uuxYmFfr3l2nxE+9e/4B/IEypcKkGTDniae2
bnGU48WQ9cGwqYi4scVWxKFArkAcGBEUs1TT4HYdXyWw4F2Vj+WGL0SY77oVuyz0tSdmxKWQU/8J
+QbQqqSyoTuyRWuOO4AjuNWkrTvf+FnBEe7x047hCUAlAhqRrtWANvcaGiPF0A+pOyHo/e+LzV1Z
qsbeyJNKtAuiCFRTdeJhNbanWZPNfo5DW9lSfengni3IVDoBlMbHfWlQT4ZFsjgvXE3rkn42VS4u
8jBoBF9uLg6ScUtpSGRziOJwFmwZ2p7zZKmtm7cTc7VizFSbPuPhC/gn1gYHsAceG+u5YpQZKAHO
VRFTrCzshkns34m1g2J751WBSX3ecbf6yvoUnwzc07b3gdhebBq6GmYSKraGA+vZFIQGunBduc0D
HjqXCzt+POPlOGIJL1Y2+W+3R2YWBNcO9KdEElf6A2yLYKPGwAKp2gLtCisnow+SRQABxkSBqanh
74uLdwYNgalVAa/9fOa2kwUR8oZXHsxqokC8bwopWlcScug6Hjj6Z6UpDxXIGp5j0X8X+1hZWuHK
SoN/XyUuPOm3tkmX9E9xTWsOJVlbwDEFWZ6vAwxDibagpcvRsE3Oz8Mx4Q9hWCd7bmIN/Osl+Rs+
nhJgMyCRGhyOWGZVPkQ3x/r/jU+PtWB0Ubwh2+6ZNC5t0lvWgP196Q7yKmzSdNMYJYLkSHt7KS8O
LNr/LOfcfYkaqVhFDbF9m5IydQfH5M1dqTPG8pPGbYFZStC+RyJy8PYbYWVYEt9MguA5VwDDkQJK
3U7Lnd6sLrIrJ/u1wG7AYdSVHYl/xPLvICKtWUEdt2pINIxgIFSQpSuYnNjCW9QB3JmXJiXmJy4A
L3+THOIeevRVy4/mVD0sRzOd1pIjfi/YaFnMFOfLFfAaw2I3GgDQnzTPhZ9doo6u7anEBI0Uo3dh
CePjmjOUgPnLSA/jz5SmPQ6WepY4fnqAQkM2F3yjqsPLxvTE3G2SSpJNP83+WWvsGolRs7cuvBly
FOX0azGDLJfdjNQdyGB/B87MXkARwnvhluMlIDXpeEpVSU+pgTddLggpXklhEbVmnHajS3DSyi88
nwPEcBsBrR81PS7D5NiXaBCefK/DDGCLBIaLIDfLozPEw1cmhRnCIuOpE2WfXfXlcEECS1sdTqPZ
AhaU9VhTCtdsfDw7RS07TkAN+LsxbzVq02VjVsgwXuBvegPlZfb/Z0XfMdsvg3NIBlHW0bv1sC/v
QBrfzTP3pMZ4SKBdq0Puo9gzb5Joo2rbvAdR3/+KLnSIgRrYcCeOEKPcyBD5QQqdBudomi20FRGQ
6fpR0jOHERbLDYPTahSYNmcL4EI/yHFi2n6J3fDVxrvH9EDJVPxwT7/Q76jrNRD58yPpIbIHUz5x
lwaPa60GUxr6WsLtLg1QbsIpOYem1iQsNJWeDJWAmiv4t6uwf3cmcIVjyf5WkkGbcsHllKdh7h/C
O0kIz9djt5LVlv/FxCCgBgeoe33AnqML56MIBax+2tveh2myO9MckOusYV434IM8XAauJLRfM+u4
NasU8tNevd1u7a2o5aJBGpGarxAbfy0vwtnyW1KcyzjDPucylQOpgOkUJvYTdxZ6hgABUSkKqz5/
YLkVF6s1QlbtRpPO2dwBmW8pu+zqb18z7Ztg+sEzRlDsQR1Ez645mGub673Bl8tl/GH0cKp7+h/p
pOu5xbSrJQ0G31WLNeZKSxdh3QmVPFi2dlF5Xj2SE0Eqs8bq3Kxc51qeYdYgpoF2BPrx4/1gO0Sz
2M533obLF2FgOMSglvUTh/60HX+ec2rDPWDzPwfLgk4Wrd208R2UoGrf96lLc6/hnQqz2CAz5rPg
Xj+4O3cUDLeK0r976LSRdufIgwQ0wV4/Rkh8f3TFTgIwJX8syZ6B9zVTq0Xgi2F22hVfpL8+m8tE
1wYJTpLxjk+jEKfBzJJpzUCQOj+7XnGGnFFrx2tPJiwg1s223dEk6PcxlcWyjsmrLc1HXq14afNg
yc1NNShAFplzue7QElrp/GtTyV96py4jET82tWRLbfy9qexGrjsj9b1nDgO4rp8Hssm2w7icYIM3
wnOpNLAJ9lg2WiOfZxbdMqAfEH6by5Tim594i3qhQKvtEB3WyVRVGE/0hrxdPADk7sA9ZMfWxYJd
p8oxWyohM3pBowwXG5bjJ76r8PXa8RmlXzC3COGiN2880gelcwcOKoen7yzC72v7r4ugrG3MzMvj
qchRKhBw9IBPnzeC5dGUfKcep2JUN348jL81VboFQ/V93GsdMvrknuko/pnPL1xUthayiHbaytV2
JZD2MaUaQ7X+whOsPViVxWgINGSJ5zHgvXJrccfkZ2Mt0Sa/Acx1J25L0P6tzcV9XQq3TJZnk2yu
zE8b4XvH4aWYgC8M5ec8QwuKa+UPXoY3IdUoTBo7Kbue6l7ELrDWeRJ+6bgEwIGD+DSq6tHywoao
c5xpP1Oyz3Goe/fRn/eTvz8al6uRXxnEVFEOxdECOItJmeVsHWzYJ54oRyjsSzhLUsB1AWANxa1Y
tkyi4urpSzLC/Q2f+DOlnqCoI4DiPsnjbIaGcBhThjLyNP+OBgN34LRzOean39Hs71skrorKY4Mj
4ZdHmfhBBrvw6Ymrar18sCYg3b3vBjIkAyxZm3qCaNbt3nNC+Lbjim2KsXzB8e+8hVt5oGX9CfzZ
otn5VZOOQAQbwFrd/fxz3Yol6cjQSCOp38MXHF6ryhoJ2VNIYLVCabDQ09ExF2UgPoCfQ0zK1THl
t2O6Eo5MIQ7urPtgPEWDQ7AC8d1n17KU1C8Qdbp0F4gvjoxgIVYY6RmDNugqtqjvI4yd2/Uvz6o8
DAGtRhKsd4XbKXP8Opb00skv2GWJ3xLWYi5Io+uhbeueJUnUvg0qKTlzUyoDVM94TxfHo10MEJgC
PnzOvOkTJD/MlOE35zKvhEA/etF6QNF/wuWYTgayntdGbFTznR2cZvZxHZomVX/vArBGumWsUqMx
/hIJlgJxSMNwiKhkdEn5QINCMpKHUZVQ9/zO313YXipsR0uVHEC1ybZz2Br0EzqRZUkGlDthLa94
/gWBBsFzOE5Yuj5eIcva5uD+71SNW9w2C6A8gWMK7YuQP9BISpHSuFgT3fw9mwEv7NaYeg1t5R30
l6ePul2k3csyQrfdk7YeuDOXdnGYJuqXYXtKctlu/I1fLsWg4ojXU4Nl0bg5hSuPBeCdFiPSf2yu
pkg5Gio2Ty26FrvZT7GeaWkkGRPz7IHIFNoCpEI5yNmXls3qhCKl2m8K3N2/EQjGn/q+KJMCyhQi
lnMC7sDXDk9GxSaVsjGOSjG6PS6QPt9xWI8hy8wU9aTzj+xgOJWZ69VIZl5LtlFha2656S0BjOV3
FTtfeH07ALgK6OZZJ267Zc7Sg8/2x9OVQZHzKo87ZJZCMOteL/wd4I+hVMxEXk+HZFv5GK7yUP0J
dyM61NBRyVUXBxPLwzlIchyYvhO0kror2dTtou3qYLFKmw92ansPk15Q91rhntq6pF5m4tr/HtZz
KYWvnekqDOOCgu8/MxRVVOVwPT7fasmbEEhaa0Yqw3leIP2WEfZFNf6od3+0p27H9vz3Pv/VtPrW
c5tBcZv0qMHpQtckK529MQ3zemdJJ7eNLZ6ruzTxwckRHybHQvfpc4la1h9M9N9aMZw42VrMrRlT
RLQuTkl5Cj9MVvaDP3xGDzaas8P1SZJC8vtI2d98nkM4TiKgTfNopRPngMBxhyRt5WwU5d0FFN5U
VFkg3psOXx25LcjGSpXiNRaZNtIv9ltJLd9iodifNwGEW9kxIqLVDsJYvYI3h8GCHXaSNaeKRFLX
iP02/RYkOZGVgmRkRaOM61Lhz+Gih5eqCP6h6turIfsskmTqDRUvY7jtsHdG604+TfylMEwxAdHM
zfClCVbR9LMmQGgr8ygTr/kpURe6JpZ4muaWaDKwP5Wg2lYGhr/Da/8lXjVr+WQFUbzgkwMEIb4g
Gdrkwu1YjGsJStvWxAKSYBp8NG7q+jioJ2rylKCEjTWcFPlgCNpYQ4yyulILCS7UQvhd3VMjXyn0
b87eNlynhUFf1Tcv7yC4wMp0UKZGt2ysE9rZ+7ef85AQaaZP0kw8dOgfcvXwlbgoJs38a0qGtEDW
vZRppyaDIaDEGeejhcmJ+D6WvBYwINFy7NL6CIP/94==
`protect end_protected
--------------------------------------------------------------------------------
--
-- File ID     : $Id: bfm_lspcie_rc.vhd 33 2021-11-16 22:43:39Z  $
-- Generated   : $LastChangedDate: 2021-11-16 23:43:39 +0100 (Tue, 16 Nov 2021) $
-- Revision    : $LastChangedRevision: 33 $
--
--------------------------------------------------------------------------------

Library IEEE;
Use IEEE.std_logic_1164.all;

Entity pcs_pipe_top is
   generic (
      g_no_scrambling   : std_logic := '0'
      );
   port(
      refclkp              : in  std_logic;         
      refclkn              : in  std_logic;         
      ffc_quad_rst         : in  std_logic := '0';     
      RESET_n              : in  std_logic;   
      pcie_ip_rstn         : out std_logic;      

      hdinp0               : in  std_logic;         
      hdinn0               : in  std_logic;         
      hdoutp0              : out std_logic;           
      hdoutn0              : out std_logic;           
      RxValid_0            : out std_logic;           
      RxElecIdle_0         : out std_logic;           
      TxData_0             : in  std_logic_vector(7 downto 0); 
      RxData_0             : out std_logic_vector(7 downto 0); 
      TxElecIdle_0         : in  std_logic; 
      TxCompliance_0       : in  std_logic; 
      TxDataK_0            : in  std_logic_vector(0 downto 0); 
      RxDataK_0            : out std_logic_vector(0 downto 0); 
      RxStatus_0           : out std_logic_vector(2 downto 0); 
      RxPolarity_0         : in  std_logic;         

      hdinp1               : in  std_logic := '0';         
      hdinn1               : in  std_logic := '0';         
      hdoutp1              : out std_logic;           
      hdoutn1              : out std_logic;           
      RxValid_1            : out std_logic;           
      RxElecIdle_1         : out std_logic;           
      TxData_1             : in  std_logic_vector(7 downto 0) := "00000000"; 
      RxData_1             : out std_logic_vector(7 downto 0); 
      TxElecIdle_1         : in  std_logic := '0'; 
      TxCompliance_1       : in  std_logic := '0'; 
      TxDataK_1            : in  std_logic_vector(0 downto 0) := "0"; 
      RxDataK_1            : out std_logic_vector(0 downto 0); 
      RxStatus_1           : out std_logic_vector(2 downto 0); 
      RxPolarity_1         : in  std_logic := '0';      

      hdinp2               : in  std_logic := '0';         
      hdinn2               : in  std_logic := '0';         
      hdoutp2              : out std_logic;           
      hdoutn2              : out std_logic;           
      RxValid_2            : out std_logic;           
      RxElecIdle_2         : out std_logic;           
      TxData_2             : in  std_logic_vector(7 downto 0):= "00000000"; 
      RxData_2             : out std_logic_vector(7 downto 0); 
      TxElecIdle_2         : in  std_logic := '0'; 
      TxCompliance_2       : in  std_logic := '0'; 
      TxDataK_2            : in  std_logic_vector(0 downto 0) := "0"; 
      RxDataK_2            : out std_logic_vector(0 downto 0); 
      RxStatus_2           : out std_logic_vector(2 downto 0); 
      RxPolarity_2         : in  std_logic := '0';      
      
      hdinp3               : in  std_logic := '0';         
      hdinn3               : in  std_logic := '0';         
      hdoutp3              : out std_logic;           
      hdoutn3              : out std_logic;           
      RxValid_3            : out std_logic;           
      RxElecIdle_3         : out std_logic;           
      TxData_3             : in  std_logic_vector(7 downto 0):= "00000000"; 
      RxData_3             : out std_logic_vector(7 downto 0); 
      TxElecIdle_3         : in  std_logic := '0'; 
      TxCompliance_3       : in  std_logic := '0'; 
      TxDataK_3            : in  std_logic_vector(0 downto 0) := "0"; 
      RxDataK_3            : out std_logic_vector(0 downto 0); 
      RxStatus_3           : out std_logic_vector(2 downto 0); 
      RxPolarity_3         : in  std_logic := '0';      
                  
      scisel_0             : in  std_logic;         
      scien_0              : in  std_logic;         
      scisel_1             : in  std_logic := '0';         
      scien_1              : in  std_logic := '0';  
      scisel_2             : in  std_logic := '0';         
      scien_2              : in  std_logic := '0';   
      scisel_3             : in  std_logic := '0';         
      scien_3              : in  std_logic := '0';                
      sciwritedata         : in  std_logic_vector(7 downto 0);
      sciaddress           : in  std_logic_vector(5 downto 0);
      scireaddata          : out std_logic_vector(7 downto 0);
      sciselaux            : in  std_logic;
      scienaux             : in  std_logic;
      scird                : in  std_logic;
      sciwstn              : in  std_logic;
      ffs_plol             : out std_logic;
      ffs_rlol_ch0         : out std_logic;

      flip_lanes           : in  std_logic := '0';                          
      PCLK                 : out std_logic;           
      PCLK_by_2            : out std_logic;           
      TxDetectRx_Loopback  : in  std_logic;         
      PhyStatus            : out std_logic;           
      PowerDown            : in  std_logic_vector(1 downto 0); 

      ctc_disable          : in  std_logic;         
      phy_ltssm_state      : in  std_logic_vector(3 downto 0) := (others => '0'); 
      phy_l0               : in  std_logic := '0';  
      phy_cfgln            : in  std_logic_vector(3 downto 0)
    );
End Entity pcs_pipe_top;
--------------------------------------------------------------------------------
--
-- File ID     : $Id: bfm_lspcie_rc.vhd 33 2021-11-16 22:43:39Z  $
-- Generated   : $LastChangedDate: 2021-11-16 23:43:39 +0100 (Tue, 16 Nov 2021) $
-- Revision    : $LastChangedRevision: 33 $
--
--------------------------------------------------------------------------------
Use WORK.bfm_lspcie_rc_types_pkg.all;

Architecture Bhv of pcs_pipe_top is
   Component bfm_lspcie_rc
      Generic (
         g_no_scrambling   : std_logic;
         g_path_root       : string;
         g_tlm_time_out    : time := 100 us;
         g_trace_label     : string := "PCIE_X1";
         g_unit_id         : natural := 1
         );
      Port (     
         i_clk_250                  : in  std_logic;
         i_rst_n                    : in std_logic;                        -- asynchronous system reset.

         i_rxp_data_0               : in  std_logic_vector(7 downto 0);
         i_rxp_data_k_0             : in  std_logic;
         i_rxp_data_1               : in  std_logic_vector(7 downto 0);
         i_rxp_data_k_1             : in  std_logic;
         i_rxp_data_2               : in  std_logic_vector(7 downto 0);
         i_rxp_data_k_2             : in  std_logic;
         i_rxp_data_3               : in  std_logic_vector(7 downto 0);
         i_rxp_data_k_3             : in  std_logic;

            -- PCIe Differential Signals
         i_refclkp                  : in  std_logic   := '0';   
         i_refclkn                  : in  std_logic   := '1';   
         i_hdinp0                   : in  std_logic   := '0';      
         i_hdinn0                   : in  std_logic   := '0'; 
         i_hdinp1                   : in  std_logic   := '0';      
         i_hdinn1                   : in  std_logic   := '0'; 
         i_hdinp2                   : in  std_logic   := '0';      
         i_hdinn2                   : in  std_logic   := '0'; 
         i_hdinp3                   : in  std_logic   := '0';      
         i_hdinn3                   : in  std_logic   := '0'; 

            -- Outputs
         o_dl_up                    : out std_logic;                       -- Data Link Layer is UP 
         o_end_sim                  : out std_logic;
         o_hdoutp0                  : out std_logic; 
         o_hdoutn0                  : out std_logic; 
         o_hdoutp1                  : out std_logic; 
         o_hdoutn1                  : out std_logic; 
         o_hdoutp2                  : out std_logic; 
         o_hdoutn2                  : out std_logic; 
         o_hdoutp3                  : out std_logic; 
         o_hdoutn3                  : out std_logic;             

         o_trc_ca_cplh              : out std_logic_vector(8 downto 0);      
         o_trc_ca_cpld              : out std_logic_vector(12 downto 0);   
         o_trc_ca_nph               : out std_logic_vector(8 downto 0);      
         o_trc_ca_npd               : out std_logic_vector(12 downto 0);     
         o_trc_ca_ph                : out std_logic_vector(8 downto 0);      
         o_trc_ca_pd                : out std_logic_vector(12 downto 0);      
         o_trc_phy_ltssm_state      : out std_logic_vector(3 downto 0);
         o_trc_phy_ltssm_substate   : out std_logic_vector(2 downto 0);
         o_trc_rx_st_vc0            : out std_logic;
         o_trc_rx_data_vc0          : out std_logic_vector(63 downto 0);
         o_trc_rx_end_vc0           : out std_logic;
         o_trc_tlp_rdy              : out std_logic;
         o_trc_tlp_req              : out std_logic;         
         o_trc_tx_st_vc0            : out std_logic;
         o_trc_tx_data_vc0          : out std_logic_vector(63 downto 0);  
         o_trc_tx_end_vc0           : out std_logic;
         o_txp_data_0               : out std_logic_vector(7 downto 0);
         o_txp_data_k_0             : out std_logic;
         o_txp_data_1               : out std_logic_vector(7 downto 0);
         o_txp_data_k_1             : out std_logic;
         o_txp_data_2               : out std_logic_vector(7 downto 0);
         o_txp_data_k_2             : out std_logic;
         o_txp_data_3               : out std_logic_vector(7 downto 0);
         o_txp_data_k_3             : out std_logic
         );
   End Component;

   Component bfm_pipe_fsm 
      Port(
         i_rst_ext_n          : in  std_logic;
         o_pcie_ip_rst_n      : out std_logic;

         i_ctl_upstream       : in  std_logic := '0';
         i_hdinn              : in  std_logic_vector;
         i_hdinp              : in  std_logic_vector;
         i_ltssm_state        : in  std_logic_vector(3 downto 0)  := (others => '0');
         i_power_down         : in  std_logic_vector(1 downto 0);
         i_rxp_data           : in  std_logic_vector(7 downto 0)  := (others => '0');
         i_rxp_data_k         : in  std_logic := '0';         
         i_stim_end_sim       : in  std_logic;
         i_txp_compliance     : in  std_logic_vector;
         i_txp_data           : in  std_logic_vector(7 downto 0)  := (others => '0');
         i_txp_data_k         : in  std_logic := '0';
         i_txp_detect_rx_lb   : in  std_logic;
         i_txp_elec_idle      : in  std_logic_vector;

         o_clk_125            : out std_logic;
         o_clk_250            : out std_logic;
         o_no_pcie_train      : out std_logic;
         o_phy_status         : out std_logic;
         o_rst_synced_n       : out std_logic;
         o_rxp_elec_idle      : out std_logic_vector;
         o_rxp_status         : out t_slv3_array;
         o_rxp_valid          : out std_logic_vector;
         o_txp_data           : out std_logic_vector(7 downto 0);
         o_txp_data_k         : out std_logic
         );
   End Component;
   

   Component pcie_scrmb
      Port (
         i_clk       : in  std_logic;
         i_rst_n     : in  std_logic;
         i_din       : in  std_logic_vector(7 downto 0);
         i_din_k     : in  std_logic;

         o_dout      : out std_logic_vector(7 downto 0);
         o_dout_k    : out std_logic
         );
   End Component;
   
   
   signal s_clk_125                    : std_logic := '0';
   signal s_clk_250                    : std_logic := '0';
   signal s_hdin_n                     : std_logic_vector(3 downto 0);
   signal s_hdin_p                     : std_logic_vector(3 downto 0);
   signal s_rst_n                      : std_logic;
   signal s_rx_data                    : std_logic_vector(31 downto 0);
   signal s_rx_data_k                  : std_logic_vector(3 downto 0);
   signal s_rxp_data_0                 : std_logic_vector(7 downto 0);
   signal s_rxp_data_1                 : std_logic_vector(7 downto 0);
   signal s_rxp_data_2                 : std_logic_vector(7 downto 0);
   signal s_rxp_data_3                 : std_logic_vector(7 downto 0);
   signal s_rxp_data_k_0               : std_logic;
   signal s_rxp_data_k_1               : std_logic;
   signal s_rxp_data_k_2               : std_logic;
   signal s_rxp_data_k_3               : std_logic;
   signal s_rxp_elec_idle              : std_logic_vector(3 downto 0);
   signal s_rxp_status                 : t_slv3_array(3 downto 0);
   signal s_rxp_valid                  : std_logic_vector(3 downto 0);
   signal s_stim_end_sim               : std_logic;  
   signal s_txp_compliance             : std_logic_vector(3 downto 0);
   signal s_txp_elec_idle              : std_logic_vector(3 downto 0);
   signal s_u1_dl_up                   : std_logic;
   signal s_u1_trc_ca_cplh             : std_logic_vector(8 downto 0);
   signal s_u1_trc_ca_cpld             : std_logic_vector(12 downto 0);
   signal s_u1_trc_ca_nph              : std_logic_vector(8 downto 0);
   signal s_u1_trc_ca_npd              : std_logic_vector(12 downto 0);
   signal s_u1_trc_ca_ph               : std_logic_vector(8 downto 0);
   signal s_u1_trc_ca_pd               : std_logic_vector(12 downto 0);
   signal s_u1_trc_phy_ltssm_state     : std_logic_vector(3 downto 0);
   signal s_u1_trc_phy_ltssm_substate  : std_logic_vector(2 downto 0);
   signal s_u1_trc_rx_st_vc0           : std_logic;
   signal s_u1_trc_rx_data_vc0         : std_logic_vector(63 downto 0);
   signal s_u1_trc_rx_end_vc0          : std_logic;
   signal s_u1_trc_tlp_rdy             : std_logic;
   signal s_u1_trc_tlp_req             : std_logic;
   signal s_u1_trc_tx_st_vc0           : std_logic;
   signal s_u1_trc_tx_data_vc0         : std_logic_vector(63 downto 0);
   signal s_u1_trc_tx_end_vc0          : std_logic;
   signal s_u3_rx_data                 : std_logic_vector(7 downto 0);
   signal s_u3_rx_data_k               : std_logic;
   signal s_u4_rx_data                 : std_logic_vector(7 downto 0);
   signal s_u4_rx_data_k               : std_logic;   
   signal s_u11_phy_status             : std_logic;
   signal s_u11_rxp_elec_idle          : std_logic_vector(3 downto 0);
   signal s_u11_rxp_valid              : std_logic_vector(3 downto 0); 
   signal s_u11_rxp_status             : t_slv3_array(3 downto 0);
    
Begin
   hdoutp0        <= '0';
   hdoutn0        <= '1';
   RxData_0       <= s_rx_data(7 downto 0) after 2ps;
   RxDataK_0(0)   <= s_rx_data_k(0) after 2ps;
   RxValid_0      <= s_u11_rxp_valid(0) after 2ps;
   RxElecIdle_0   <= s_u11_rxp_elec_idle(0) after 2ps;
   RxStatus_0     <= s_u11_rxp_status(0) after 2ps;

   hdoutp1        <= '0';
   hdoutn1        <= '1';
   RxData_1       <= s_rx_data(15 downto 8) after 2ps;
   RxDataK_1(0)   <= s_rx_data_k(1) after 2ps;
   RxValid_1      <= s_u11_rxp_valid(1) after 2ps;
   RxElecIdle_1   <= s_u11_rxp_elec_idle(1) after 2ps;
   RxStatus_1     <= s_u11_rxp_status(1) after 2ps;
   
   hdoutp2        <= '0';
   hdoutn2        <= '1';
   RxData_2       <= s_rx_data(23 downto 16) after 2ps;
   RxDataK_2(0)   <= s_rx_data_k(2) after 2ps;
   RxValid_2      <= s_u11_rxp_valid(2) after 2ps;
   RxElecIdle_2   <= s_u11_rxp_elec_idle(2) after 2ps;
   RxStatus_2     <= s_u11_rxp_status(2) after 2ps;   
      
   hdoutp3        <= '0';
   hdoutn3        <= '1';
   RxData_3       <= s_rx_data(31 downto 24) after 2ps;
   RxDataK_3(0)   <= s_rx_data_k(3) after 2ps;
   RxValid_3      <= s_u11_rxp_valid(3) after 2ps;
   RxElecIdle_3   <= s_u11_rxp_elec_idle(3) after 2ps;
   RxStatus_3     <= s_u11_rxp_status(3) after 2ps;
         
   scireaddata    <= (others => '0');
   ffs_plol       <= '0';
   ffs_rlol_ch0   <= '0';
   PCLK           <= s_clk_250;
   PCLK_by_2      <= s_clk_125 after 1 ps;
   PhyStatus      <= s_u11_phy_status after 2ps;
   
   --s_hdin_n          <= (others => '0');
   --s_hdin_p          <= (0 => '1', others => '0');
   s_hdin_n          <= hdinn3 & hdinn2 & hdinn1 & hdinn0;
   s_hdin_p          <= hdinp3 & hdinp2 & hdinp1 & hdinp0;   
   s_txp_compliance  <= TxCompliance_3 & TxCompliance_2 & TxCompliance_1 & TxCompliance_0;
   s_txp_elec_idle(3)   <= '1' when TxElecIdle_3 = '1' else '0';
   s_txp_elec_idle(2)   <= '1' when TxElecIdle_2 = '1' else '0';
   s_txp_elec_idle(1)   <= '1' when TxElecIdle_1 = '1' else '0';
   s_txp_elec_idle(0)   <= '1' when TxElecIdle_0 = '1' else '0';

   s_rxp_data_0      <= TxData_0 after 1ps;
   s_rxp_data_k_0    <= TxDataK_0(0) after 1ps;
   s_rxp_data_1      <= TxData_1 after 100ps;
   s_rxp_data_k_1    <= TxDataK_1(0) after 1ps;
   s_rxp_data_2      <= TxData_2 after 1ps;
   s_rxp_data_k_2    <= TxDataK_2(0) after 1ps;
   s_rxp_data_3      <= TxData_3 after 1ps;
   s_rxp_data_k_3    <= TxDataK_3(0) after 1ps;
   
      --    ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   U1_BFM: bfm_lspcie_rc
      Generic Map (
         g_no_scrambling   => g_no_scrambling,
         g_path_root       => Bhv'path_name
         )
      Port Map (
         i_clk_250                  => s_clk_250,
         i_rst_n                    => RESET_n,
         i_hdinp0                   => hdinp0,
         i_hdinn0                   => hdinn0,
         i_hdinp1                   => hdinp1,
         i_hdinn1                   => hdinn1,
         i_hdinp2                   => hdinp2,
         i_hdinn2                   => hdinn2,
         i_hdinp3                   => hdinp3,
         i_hdinn3                   => hdinn3,    
         i_rxp_data_0               => s_rxp_data_0, 
         i_rxp_data_k_0             => s_rxp_data_k_0,
         i_rxp_data_1               => s_rxp_data_1,  
         i_rxp_data_k_1             => s_rxp_data_k_1,
         i_rxp_data_2               => s_rxp_data_2,  
         i_rxp_data_k_2             => s_rxp_data_k_2,
         i_rxp_data_3               => s_rxp_data_3,  
         i_rxp_data_k_3             => s_rxp_data_k_3,
                           
         o_dl_up                    => s_u1_dl_up,
         o_end_sim                  => s_stim_end_sim,
         o_trc_ca_cplh              => s_u1_trc_ca_cplh,
         o_trc_ca_cpld              => s_u1_trc_ca_cpld,
         o_trc_ca_nph               => s_u1_trc_ca_nph,
         o_trc_ca_npd               => s_u1_trc_ca_npd,
         o_trc_ca_ph                => s_u1_trc_ca_ph,
         o_trc_ca_pd                => s_u1_trc_ca_pd,
         o_trc_phy_ltssm_state      => s_u1_trc_phy_ltssm_state,
         o_trc_phy_ltssm_substate   => s_u1_trc_phy_ltssm_substate,
         o_trc_rx_st_vc0            => s_u1_trc_rx_st_vc0,
         o_trc_rx_data_vc0          => s_u1_trc_rx_data_vc0,
         o_trc_rx_end_vc0           => s_u1_trc_rx_end_vc0,
         o_trc_tlp_rdy              => s_u1_trc_tlp_rdy,
         o_trc_tlp_req              => s_u1_trc_tlp_req,
         o_trc_tx_st_vc0            => s_u1_trc_tx_st_vc0,
         o_trc_tx_data_vc0          => s_u1_trc_tx_data_vc0,
         o_trc_tx_end_vc0           => s_u1_trc_tx_end_vc0,
         o_txp_data_0               => s_rx_data(7 downto 0),
         o_txp_data_k_0             => s_rx_data_k(0),
         o_txp_data_1               => s_rx_data(15 downto 8),
         o_txp_data_k_1             => s_rx_data_k(1),
         o_txp_data_2               => s_rx_data(23 downto 16),
         o_txp_data_k_2             => s_rx_data_k(2),
         o_txp_data_3               => s_rx_data(31 downto 24),
         o_txp_data_k_3             => s_rx_data_k(3)                  
         );
         

   U2_PIPE:
      -- This is the PIPE interface for the DUT
   bfm_pipe_fsm 
      Port Map (
         i_rst_ext_n          => RESET_n,
         o_pcie_ip_rst_n      => pcie_ip_rstn,

         i_hdinn              => s_hdin_n,
         i_hdinp              => s_hdin_p,
         i_power_down         => PowerDown,
         i_rxp_data           => s_rx_data(7 downto 0),
         i_rxp_data_k         => s_rx_data_k(0),           
         i_stim_end_sim       => s_stim_end_sim,
         i_txp_compliance     => s_txp_compliance,
         i_txp_detect_rx_lb   => TxDetectRx_Loopback,
         i_txp_elec_idle      => s_txp_elec_idle,

         o_clk_125            => s_clk_125,
         o_clk_250            => s_clk_250,
         o_rst_synced_n       => s_rst_n,
         o_no_pcie_train      => open,
         o_phy_status         => s_u11_phy_status,
         o_rxp_elec_idle      => s_u11_rxp_elec_idle,
         o_rxp_status         => s_u11_rxp_status,
         o_rxp_valid          => s_u11_rxp_valid
         );
         
   U3_RX_SCRMB:
   pcie_scrmb
      Port Map(
         i_clk       => s_clk_250,
         i_rst_n     => RESET_n,
         i_din       => s_rx_data(7 downto 0),
         i_din_k     => s_rx_data_k(0),

         o_dout      => s_u3_rx_data,
         o_dout_k    => s_u3_rx_data_k
         );
         
   U4_TX_SCRMB:
   pcie_scrmb
      Port Map(
         i_clk       => s_clk_250,
         i_rst_n     => RESET_n,
         i_din       => s_rxp_data_0,
         i_din_k     => s_rxp_data_k_0,

         o_dout      => s_u4_rx_data,
         o_dout_k    => s_u4_rx_data_k
         );         
End Bhv;

--
--------------------------------------------------------------------------------
--
-- File ID     : $Id: bfm_lspcie_rc.vhd 33 2021-11-16 22:43:39Z  $
-- Generated   : $LastChangedDate: 2021-11-16 23:43:39 +0100 (Tue, 16 Nov 2021) $
-- Revision    : $LastChangedRevision: 33 $
--
--------------------------------------------------------------------------------
Library IEEE;
Use IEEE.std_logic_1164.all;
Use WORK.bfm_lspcie_rc_constants_pkg.all;
Use WORK.bfm_lspcie_rc_tlm_lib_pkg.all;
Use WORK.bfm_lspcie_rc_types_pkg.all;
Use WORK.bfm_random_data_pkg.all;

Package pcie_vhdl_test_case_pkg is
   procedure run_test(signal clk       : in    std_logic;
                      signal sv        : inout t_bfm_stim;
                      signal rv        : in    t_bfm_resp;
                             id        : in    natural := 0); 

End pcie_vhdl_test_case_pkg;
--
--------------------------------------------------------------------------------
--
-- File ID     : $Id: bfm_lspcie_rc.vhd 33 2021-11-16 22:43:39Z  $
-- Generated   : $LastChangedDate: 2021-11-16 23:43:39 +0100 (Tue, 16 Nov 2021) $
-- Revision    : $LastChangedRevision: 33 $
--
--------------------------------------------------------------------------------

Library IEEE;

Use IEEE.std_logic_1164.all;
Use STD.env.all;
Use STD.textio.all;
Use WORK.bfm_lspcie_rc_tlm_lib_pkg.all;
Use WORK.bfm_lspcie_rc_utils_pkg.all;
Use WORK.bfm_lspcie_rc_types_pkg.all;

Entity pcie_stim_vhdl is
   Generic (
      g_path_root          : string
      );
   Port (
      i_clk_125            : in  std_logic;
      i_rst_n              : in  std_logic;
     
      i_bfm_resp           : in  t_bfm_resp;
      i_dl_up              : in  std_logic;
      
      o_bfm_stim           : inout t_bfm_stim := c_bfm_stim_init
      );
End pcie_stim_vhdl;

--
--------------------------------------------------------------------------------
--
-- File ID     : $Id: bfm_lspcie_rc.vhd 33 2021-11-16 22:43:39Z  $
-- Generated   : $LastChangedDate: 2021-11-16 23:43:39 +0100 (Tue, 16 Nov 2021) $
-- Revision    : $LastChangedRevision: 33 $
--
--------------------------------------------------------------------------------
--    To interact with other BFMs or for more complex verification scenarios
--    for instance, the user can modify this file
--
--    Normally, this file just calls the test-case through the 'run_test' call
--    below.
--------------------------------------------------------------------------------

Use WORK.pcie_vhdl_test_case_pkg.all;

Architecture Bhv of pcie_stim_vhdl is

Begin

   R_MAIN:
   process
      variable v_line   : line;
   begin      
      wait for 0 ns;
      wait until (i_rst_n = '1');
      idle(i_clk_125, 8);
         
      wait until (i_dl_up = '1');
      idle(i_clk_125);
      msgd_set_slot_power_limit(i_clk_125, o_bfm_stim, i_bfm_resp, value => X"02", scale => "01");

         -- Call the Test Case
      run_test(i_clk_125, o_bfm_stim, i_bfm_resp); 

      idle(i_clk_125, 128);
      
      assert false report LF & LF & "        +++ Game Over +++" & LF & LF severity note;             
      wait for 5 ns;
      stop(0);
   end process;   

End Bhv;

--
--------------------------------------------------------------------------------
--
-- File ID     : $Id: bfm_lspcie_rc.vhd 33 2021-11-16 22:43:39Z  $
-- Generated   : $LastChangedDate: 2021-11-16 23:43:39 +0100 (Tue, 16 Nov 2021) $
-- Revision    : $LastChangedRevision: 33 $
--
--------------------------------------------------------------------------------

Package Body pcie_vhdl_test_case_pkg is
   procedure run_test(signal clk : in    std_logic;
                      signal sv  : inout t_bfm_stim;
                      signal rv  : in    t_bfm_resp;
                             id  : in    natural := 0) is
   begin
      wait;
   end procedure; 

End pcie_vhdl_test_case_pkg;
