Entity versa_ecp5_tb is
End versa_ecp5_tb;
