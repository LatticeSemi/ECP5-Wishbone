
--
--------------------------------------------------------------------------------
--
-- File ID     : $Id: pcie_vhdl_test_case-pb.vhd 33 2021-11-16 22:43:39Z  $
-- Generated   : $LastChangedDate: 2021-11-16 23:43:39 +0100 (Tue, 16 Nov 2021) $
-- Revision    : $LastChangedRevision: 33 $
--
--------------------------------------------------------------------------------

Package Body pcie_vhdl_test_case_pkg is
   procedure run_test(signal clk : in    std_logic;
                      signal sv  : inout t_bfm_stim;
                      signal rv  : in    t_bfm_resp;
                             id  : in    natural := 0) is
   begin
      wait;
   end procedure; 

End pcie_vhdl_test_case_pkg;
