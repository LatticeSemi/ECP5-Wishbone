`timescale 1ns / 1 ps
module pcie_vlog_test_case;
`include "bfm_lspcie_rc_tlm_lib.v"
 
      integer v_reg_val;
   initial begin
      #1;
      end
endmodule
