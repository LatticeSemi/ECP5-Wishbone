
--    
--    Copyright Ingenieurbuero Gardiner, 2021
--       https://www.ib-gardiner.eu
--       techsupport@ib-gardiner.eu
--
--    All Rights Reserved
--   
--------------------------------------------------------------------------------
--
-- File ID    : $Id: lscc_pcie_x1_ip-a_rtl.vhd 46 2021-11-18 22:45:40Z  $
-- Generated  : $LastChangedDate: 2021-11-18 23:45:40 +0100 (Thu, 18 Nov 2021) $
-- Revision   : $LastChangedRevision: 46 $
--
--------------------------------------------------------------------------------
--
-- Description : 
--
--------------------------------------------------------------------------------
Use WORK.tspc_utils.all;

Architecture Rtl of lscc_pcie_x1_ip is
   signal s_rtl_inta_n              : std_logic;
 --signal s_u1_refclk               : std_logic;
   signal s_u2_rst_n                : std_logic;

   Component tspc_rst_gen_yog4
      Generic (
         g_rst_count    : positive := 16#9C4#
         );
      Port (
         i_clk       : in  std_logic;
         i_trip_ev   : in  std_logic;
         
         o_rst_n     : out std_logic
         );
   End Component;

   Component pcie_x1_e5
         -- Module generated by Clarity. Component name must match Clarity name
         --
         -- Assumption : instance name of PCIe core is x_pcie
         --              instance name of ref clock is x_cref
         -- If these are different the port-names below must be updated accordingly
         -- or the ports on the clarity design renamed.
         -- 
         -- Otherwise, there is normally no need to change the port declarations
      Port (
         x_cref_refclkn                : in  std_logic;
         x_cref_refclkp                : in  std_logic;
         x_pcie_cmpln_tout             : in  std_logic;
         x_pcie_cmpltr_abort_np        : in  std_logic;
         x_pcie_cmpltr_abort_p         : in  std_logic;
         x_pcie_flip_lanes             : in  std_logic;
         x_pcie_force_disable_scr      : in  std_logic;
         x_pcie_force_lsm_active       : in  std_logic;
         x_pcie_force_phy_status       : in  std_logic;
         x_pcie_force_rec_ei           : in  std_logic;
         x_pcie_hdinn0                 : in  std_logic;
         x_pcie_hdinp0                 : in  std_logic;
         x_pcie_hl_disable_scr         : in  std_logic;
         x_pcie_hl_gto_cfg             : in  std_logic;
         x_pcie_hl_gto_det             : in  std_logic;
         x_pcie_hl_gto_dis             : in  std_logic;
         x_pcie_hl_gto_hrst            : in  std_logic;
         x_pcie_hl_gto_l0stx           : in  std_logic;
         x_pcie_hl_gto_l0stxfts        : in  std_logic;
         x_pcie_hl_gto_l1              : in  std_logic;
         x_pcie_hl_gto_l2              : in  std_logic;
         x_pcie_hl_gto_lbk             : in  std_logic;
         x_pcie_hl_gto_rcvry           : in  std_logic;
         x_pcie_hl_snd_beacon          : in  std_logic;
         x_pcie_inta_n                 : in  std_logic;
         x_pcie_msi                    : in  std_logic_vector(7 downto 0);
         x_pcie_no_pcie_train          : in  std_logic;
         x_pcie_np_req_pend            : in  std_logic;
         x_pcie_npd_buf_status_vc0     : in  std_logic;
         x_pcie_npd_num_vc0            : in  std_logic_vector(7 downto 0);
         x_pcie_npd_processed_vc0      : in  std_logic;
         x_pcie_nph_buf_status_vc0     : in  std_logic;
         x_pcie_nph_processed_vc0      : in  std_logic;
         x_pcie_pd_buf_status_vc0      : in  std_logic;
         x_pcie_pd_num_vc0             : in  std_logic_vector(7 downto 0);
         x_pcie_pd_processed_vc0       : in  std_logic;
         x_pcie_ph_buf_status_vc0      : in  std_logic;
         x_pcie_ph_processed_vc0       : in  std_logic;
         x_pcie_pll_refclki            : in  std_logic;
         x_pcie_pme_status             : in  std_logic;
         x_pcie_rst_n                  : in  std_logic;
         x_pcie_rxrefclk               : in  std_logic;
         x_pcie_sci_addr               : in  std_logic_vector(5 downto 0);
         x_pcie_sci_en                 : in  std_logic;
         x_pcie_sci_en_dual            : in  std_logic;
         x_pcie_sci_rd                 : in  std_logic;
         x_pcie_sci_sel                : in  std_logic;
         x_pcie_sci_sel_dual           : in  std_logic;
         x_pcie_sci_wrdata             : in  std_logic_vector(7 downto 0);
         x_pcie_sci_wrn                : in  std_logic;
         x_pcie_tx_data_vc0            : in  std_logic_vector(15 downto 0);
         x_pcie_tx_dllp_val            : in  std_logic_vector(1 downto 0);
         x_pcie_tx_end_vc0             : in  std_logic;
         x_pcie_tx_lbk_data            : in  std_logic_vector(15 downto 0);
         x_pcie_tx_lbk_kcntl           : in  std_logic_vector(1 downto 0);
         x_pcie_tx_nlfy_vc0            : in  std_logic;
         x_pcie_tx_pmtype              : in  std_logic_vector(2 downto 0);
         x_pcie_tx_req_vc0             : in  std_logic;
         x_pcie_tx_st_vc0              : in  std_logic;
         x_pcie_tx_vsd_data            : in  std_logic_vector(23 downto 0);
         x_pcie_unexp_cmpln            : in  std_logic;
         x_pcie_ur_np_ext              : in  std_logic;
         x_pcie_ur_p_ext               : in  std_logic;

         x_cref_refclko                : out std_logic;
         x_pcie_bus_num                : out std_logic_vector(7 downto 0);
         x_pcie_cmd_reg_out            : out std_logic_vector(5 downto 0);
         x_pcie_dev_cntl_out           : out std_logic_vector(14 downto 0);
         x_pcie_dev_num                : out std_logic_vector(4 downto 0);
         x_pcie_dl_active              : out std_logic;
         x_pcie_dl_inactive            : out std_logic;
         x_pcie_dl_init                : out std_logic;
         x_pcie_dl_up                  : out std_logic;
         x_pcie_func_num               : out std_logic_vector(2 downto 0);
         x_pcie_hdoutn0                : out std_logic;
         x_pcie_hdoutp0                : out std_logic;
         x_pcie_lnk_cntl_out           : out std_logic_vector(7 downto 0);
         x_pcie_mm_enable              : out std_logic_vector(2 downto 0);
         x_pcie_msi_enable             : out std_logic;
         x_pcie_phy_ltssm_state        : out std_logic_vector(3 downto 0);
         x_pcie_phy_pol_compliance     : out std_logic;
         x_pcie_pm_power_state         : out std_logic_vector(1 downto 0);
         x_pcie_pme_en                 : out std_logic;
         x_pcie_rx_bar_hit             : out std_logic_vector(6 downto 0);
         x_pcie_rx_data_vc0            : out std_logic_vector(15 downto 0);
         x_pcie_rx_end_vc0             : out std_logic;
         x_pcie_rx_lbk_data            : out std_logic_vector(15 downto 0);
         x_pcie_rx_lbk_kcntl           : out std_logic_vector(1 downto 0);
         x_pcie_rx_malf_tlp_vc0        : out std_logic;
         x_pcie_rx_st_vc0              : out std_logic;
         x_pcie_rx_us_req_vc0          : out std_logic;
         x_pcie_rxdp_dllp_val          : out std_logic_vector(1 downto 0);
         x_pcie_rxdp_pmd_type          : out std_logic_vector(2 downto 0);
         x_pcie_rxdp_vsd_data          : out std_logic_vector(23 downto 0);
         x_pcie_sci_int                : out std_logic;
         x_pcie_sci_rddata             : out std_logic_vector(7 downto 0);
         x_pcie_serdes_pdb             : out std_logic;
         x_pcie_serdes_rst_dual_c      : out std_logic;
         x_pcie_sys_clk_125            : out std_logic;
         x_pcie_tx_ca_cpl_recheck_vc0  : out std_logic;
         x_pcie_tx_ca_cpld_vc0         : out std_logic_vector(12 downto 0);
         x_pcie_tx_ca_cplh_vc0         : out std_logic_vector(8 downto 0);
         x_pcie_tx_ca_npd_vc0          : out std_logic_vector(12 downto 0);
         x_pcie_tx_ca_nph_vc0          : out std_logic_vector(8 downto 0);
         x_pcie_tx_ca_p_recheck_vc0    : out std_logic;
         x_pcie_tx_ca_pd_vc0           : out std_logic_vector(12 downto 0);
         x_pcie_tx_ca_ph_vc0           : out std_logic_vector(8 downto 0);
         x_pcie_tx_dllp_sent           : out std_logic;
         x_pcie_tx_lbk_rdy             : out std_logic;
         x_pcie_tx_pwrup_c             : out std_logic;
         x_pcie_tx_rdy_vc0             : out std_logic;
         x_pcie_tx_serdes_rst_c        : out std_logic
         );
   End Component;

   
   Component pcie_x1_e5g2
         -- Module generated by Clarity. Component name must match Clarity name
         --
         -- Assumption : instance name of PCIe core is x_pcie
         --              instance name of ref clock is x_cref
         -- If these are different the port-names below must be updated accordingly
         -- or the ports on the clarity design renamed.
         -- 
         -- Otherwise, there is normally no need to change the port declarations
      Port (
         x_cref_refclkn                : in  std_logic;
         x_cref_refclkp                : in  std_logic;
         x_pcie_cmpln_tout             : in  std_logic;
         x_pcie_cmpltr_abort_np        : in  std_logic;
         x_pcie_cmpltr_abort_p         : in  std_logic;
         x_pcie_flip_lanes             : in  std_logic;
         x_pcie_flr_rdy_in             : in  std_logic;
         x_pcie_force_disable_scr      : in  std_logic;
         x_pcie_force_lsm_active       : in  std_logic;
         x_pcie_force_phy_status       : in  std_logic;
         x_pcie_force_rec_ei           : in  std_logic;
         x_pcie_hdinn0                 : in  std_logic;
         x_pcie_hdinp0                 : in  std_logic;
         x_pcie_hl_disable_scr         : in  std_logic;
         x_pcie_hl_gto_cfg             : in  std_logic;
         x_pcie_hl_gto_det             : in  std_logic;
         x_pcie_hl_gto_dis             : in  std_logic;
         x_pcie_hl_gto_hrst            : in  std_logic;
         x_pcie_hl_gto_l0stx           : in  std_logic;
         x_pcie_hl_gto_l0stxfts        : in  std_logic;
         x_pcie_hl_gto_l1              : in  std_logic;
         x_pcie_hl_gto_l2              : in  std_logic;
         x_pcie_hl_gto_lbk             : in  std_logic_vector(1 downto 0);
         x_pcie_hl_gto_rcvry           : in  std_logic;
         x_pcie_hl_snd_beacon          : in  std_logic;
         x_pcie_inta_n                 : in  std_logic;
         x_pcie_msi                    : in  std_logic_vector(7 downto 0);
         x_pcie_no_pcie_train          : in  std_logic;
         x_pcie_np_req_pend            : in  std_logic;
         x_pcie_npd_buf_status_vc0     : in  std_logic;
         x_pcie_npd_num_vc0            : in  std_logic_vector(7 downto 0);
         x_pcie_npd_processed_vc0      : in  std_logic;
         x_pcie_nph_buf_status_vc0     : in  std_logic;
         x_pcie_nph_processed_vc0      : in  std_logic;
         x_pcie_pd_buf_status_vc0      : in  std_logic;
         x_pcie_pd_num_vc0             : in  std_logic_vector(7 downto 0);
         x_pcie_pd_processed_vc0       : in  std_logic;
         x_pcie_ph_buf_status_vc0      : in  std_logic;
         x_pcie_ph_processed_vc0       : in  std_logic;
         x_pcie_pll_refclki            : in  std_logic;
         x_pcie_pme_status             : in  std_logic;
         x_pcie_rst_n                  : in  std_logic;
         x_pcie_rxrefclk               : in  std_logic;
         x_pcie_tx_data_vc0            : in  std_logic_vector(63 downto 0);
         x_pcie_tx_dllp_val            : in  std_logic_vector(1 downto 0);
         x_pcie_tx_dwen_vc0            : in  std_logic;
         x_pcie_tx_end_vc0             : in  std_logic;
         x_pcie_tx_lbk_data            : in  std_logic_vector(63 downto 0);
         x_pcie_tx_lbk_kcntl           : in  std_logic_vector(7 downto 0);
         x_pcie_tx_nlfy_vc0            : in  std_logic;
         x_pcie_tx_pmtype              : in  std_logic_vector(2 downto 0);
         x_pcie_tx_req_vc0             : in  std_logic;
         x_pcie_tx_st_vc0              : in  std_logic;
         x_pcie_tx_vsd_data            : in  std_logic_vector(23 downto 0);
         x_pcie_unexp_cmpln            : in  std_logic;
         x_pcie_ur_np_ext              : in  std_logic;
         x_pcie_ur_p_ext               : in  std_logic;
         
         x_cref_refclko                : out std_logic;
         x_pcie_bus_num                : out std_logic_vector(7 downto 0);
         x_pcie_cmd_reg_out            : out std_logic_vector(5 downto 0);
         x_pcie_dev_cntl_2_out         : out std_logic_vector(4 downto 0);
         x_pcie_dev_cntl_out           : out std_logic_vector(14 downto 0);
         x_pcie_dev_num                : out std_logic_vector(4 downto 0);
         x_pcie_dl_active              : out std_logic;
         x_pcie_dl_inactive            : out std_logic;
         x_pcie_dl_init                : out std_logic;
         x_pcie_dl_up                  : out std_logic;
         x_pcie_func_num               : out std_logic_vector(2 downto 0);
         x_pcie_hdoutn0                : out std_logic;
         x_pcie_hdoutp0                : out std_logic;
         x_pcie_initiate_flr           : out std_logic;
         x_pcie_lnk_cntl_out           : out std_logic_vector(7 downto 0);
         x_pcie_mm_enable              : out std_logic_vector(2 downto 0);
         x_pcie_msi_enable             : out std_logic;
         x_pcie_phy_cfgln              : out std_logic_vector(1 downto 0);
         x_pcie_phy_cfgln_sum          : out std_logic_vector(2 downto 0);
         x_pcie_phy_ltssm_state        : out std_logic_vector(3 downto 0);
         x_pcie_phy_pol_compliance     : out std_logic;
         x_pcie_pm_power_state         : out std_logic_vector(1 downto 0);
         x_pcie_pme_en                 : out std_logic;
         x_pcie_rx_bar_hit             : out std_logic_vector(6 downto 0);
         x_pcie_rx_data_vc0            : out std_logic_vector(63 downto 0);
         x_pcie_rx_dwen_vc0            : out std_logic;
         x_pcie_rx_end_vc0             : out std_logic;
         x_pcie_rx_lbk_data            : out std_logic_vector(63 downto 0);
         x_pcie_rx_lbk_kcntl           : out std_logic_vector(7 downto 0);
         x_pcie_rx_malf_tlp_vc0        : out std_logic;
         x_pcie_rx_st_vc0              : out std_logic;
         x_pcie_rx_us_req_vc0          : out std_logic;
         x_pcie_rxdp_dllp_val          : out std_logic_vector(1 downto 0);
         x_pcie_rxdp_pmd_type          : out std_logic_vector(2 downto 0);
         x_pcie_rxdp_vsd_data          : out std_logic_vector(23 downto 0);
         x_pcie_sys_clk_125            : out std_logic;
         x_pcie_tx_ca_cpl_recheck_vc0  : out std_logic;
         x_pcie_tx_ca_cpld_vc0         : out std_logic_vector(12 downto 0);
         x_pcie_tx_ca_cplh_vc0         : out std_logic_vector(8 downto 0);
         x_pcie_tx_ca_npd_vc0          : out std_logic_vector(12 downto 0);
         x_pcie_tx_ca_nph_vc0          : out std_logic_vector(8 downto 0);
         x_pcie_tx_ca_p_recheck_vc0    : out std_logic;
         x_pcie_tx_ca_pd_vc0           : out std_logic_vector(12 downto 0);
         x_pcie_tx_ca_ph_vc0           : out std_logic_vector(8 downto 0);
         x_pcie_tx_dllp_sent           : out std_logic;
         x_pcie_tx_lbk_rdy             : out std_logic;
         x_pcie_tx_rdy_vc0             : out std_logic;
         x_pcie_tx_val                 : out std_logic
         );
   End Component;
   

Begin
   s_rtl_inta_n      <= not ix_int_req;

   U1_ECP3:
   if g_tech_lib = "ECP3" or g_tech_lib = "ECP2M" Generate
   
      U1_V6_X :
      if g_ip_rev_id = "V6_x" Generate   
         Component pcie_x1_ipx
               -- Module generated by ipExpress. Component name must match ipExpress name
               -- There is normally no need to change the port declarations
               
               -- References file generated by IPexpress in IP directory 
            Port (
               refclkp                 : in std_logic;
               refclkn                 : in std_logic;
               rst_n                   : in std_logic;
               flip_lanes              : in std_logic;
               hdinp0                  : in std_logic;
               hdinn0                  : in std_logic;
               hdoutp0                 : out std_logic;
               hdoutn0                 : out std_logic;
               inta_n                  : in std_logic;
               msi                     : in std_logic_vector(7 downto 0);
               force_lsm_active        : in std_logic;
               force_rec_ei            : in std_logic;
               force_phy_status        : in std_logic;
               force_disable_scr       : in std_logic;
               hl_snd_beacon           : in std_logic;
               hl_disable_scr          : in std_logic;
               hl_gto_dis              : in std_logic;
               hl_gto_det              : in std_logic;
               hl_gto_hrst             : in std_logic;
               hl_gto_l0stx            : in std_logic;
               hl_gto_l1               : in std_logic;
               hl_gto_l2               : in std_logic;
               hl_gto_l0stxfts         : in std_logic;
               hl_gto_lbk              : in std_logic;
               hl_gto_rcvry            : in std_logic;
               hl_gto_cfg              : in std_logic;
               no_pcie_train           : in std_logic;
               tx_dllp_val             : in std_logic_vector(1 downto 0);
               tx_pmtype               : in std_logic_vector(2 downto 0);
               tx_vsd_data             : in std_logic_vector(23 downto 0);
               tx_req_vc0              : in std_logic;
               tx_data_vc0             : in std_logic_vector(15 downto 0);
               tx_st_vc0               : in std_logic;
               tx_end_vc0              : in std_logic;
               tx_nlfy_vc0             : in std_logic;
               ph_buf_status_vc0       : in std_logic;
               pd_buf_status_vc0       : in std_logic;
               nph_buf_status_vc0      : in std_logic;
               npd_buf_status_vc0      : in std_logic;
               ph_processed_vc0        : in std_logic;
               pd_processed_vc0        : in std_logic;
               nph_processed_vc0       : in std_logic;
               npd_processed_vc0       : in std_logic;
               pd_num_vc0              : in std_logic_vector(7 downto 0);
               npd_num_vc0             : in std_logic_vector(7 downto 0);
               cmpln_tout              : in std_logic;
               cmpltr_abort_np         : in std_logic;
               cmpltr_abort_p          : in std_logic;
               unexp_cmpln             : in std_logic;
               ur_np_ext               : in std_logic;
               ur_p_ext                : in std_logic;
               np_req_pend             : in std_logic;
               pme_status              : in std_logic;
               tx_lbk_data             : in std_logic_vector(15 downto 0);
               tx_lbk_kcntl            : in std_logic_vector(1 downto 0);
               
               tx_lbk_rdy              : out std_logic;
               rx_lbk_data             : out std_logic_vector(15 downto 0);
               rx_lbk_kcntl            : out std_logic_vector(1 downto 0);
               tx_dllp_sent            : out std_logic;
               rxdp_pmd_type           : out std_logic_vector(2 downto 0);
               rxdp_vsd_data           : out std_logic_vector(23 downto 0);
               rxdp_dllp_val           : out std_logic_vector(1 downto 0);
               phy_pol_compliance      : out std_logic;
               phy_ltssm_state         : out std_logic_vector(3 downto 0);
               tx_rdy_vc0              : out std_logic;
               tx_ca_ph_vc0            : out std_logic_vector(8 downto 0);
               tx_ca_pd_vc0            : out std_logic_vector(12 downto 0);
               tx_ca_nph_vc0           : out std_logic_vector(8 downto 0);
               tx_ca_npd_vc0           : out std_logic_vector(12 downto 0);
               tx_ca_cplh_vc0          : out std_logic_vector(8 downto 0);
               tx_ca_cpld_vc0          : out std_logic_vector(12 downto 0);
               tx_ca_p_recheck_vc0     : out std_logic;
               tx_ca_cpl_recheck_vc0   : out std_logic;
               rx_data_vc0             : out std_logic_vector(15 downto 0);
               rx_st_vc0               : out std_logic;
               rx_end_vc0              : out std_logic;
               rx_us_req_vc0           : out std_logic;
               rx_malf_tlp_vc0         : out std_logic;
               rx_bar_hit              : out std_logic_vector(6 downto 0);
               mm_enable               : out std_logic_vector(2 downto 0);
               msi_enable              : out std_logic;
               bus_num                 : out std_logic_vector(7 downto 0);
               dev_num                 : out std_logic_vector(4 downto 0);
               func_num                : out std_logic_vector(2 downto 0);
               pm_power_state          : out std_logic_vector(1 downto 0);
               pme_en                  : out std_logic;
               cmd_reg_out             : out std_logic_vector(5 downto 0);
               dev_cntl_out            : out std_logic_vector(14 downto 0);
               lnk_cntl_out            : out std_logic_vector(7 downto 0);
               dl_inactive             : out std_logic;
               dl_init                 : out std_logic;
               dl_active               : out std_logic;
               dl_up                   : out std_logic;
               sys_clk_125             : out std_logic;
               sci_wrdata              : in std_logic_vector(7 downto 0);
               sci_addr                : in std_logic_vector(5 downto 0);
               sci_wrn                 : in std_logic;
               sci_en                  : in std_logic;
               sci_sel                 : in std_logic;
               sci_en_ch0              : in std_logic;
               sci_sel_ch0             : in std_logic;
               sci_rd                  : in std_logic;
               sci_rddata              : out std_logic_vector(7 downto 0)
               );
         End Component;      
      Begin   
         U1_PCIE:
         pcie_x1_ipx
            Port Map (
               refclkp                 => ix_refclkp,
               refclkn                 => ix_refclkn,
               rst_n                   => ix_rst_n,
               flip_lanes              => c_tie_low,
               hdinp0                  => ix_hdinp0,
               hdinn0                  => ix_hdinn0,
               hdoutp0                 => ox_hdoutp0,
               hdoutn0                 => ox_hdoutn0,
               inta_n                  => s_rtl_inta_n,
               msi                     => ix_msi_req,
               force_lsm_active        => c_tie_low,
               force_rec_ei            => c_tie_low,
               force_phy_status        => c_tie_low,
               force_disable_scr       => c_tie_low,
               hl_snd_beacon           => c_tie_low,
               hl_disable_scr          => c_tie_low,
               hl_gto_dis              => c_tie_low,
               hl_gto_det              => c_tie_low,
               hl_gto_hrst             => c_tie_low,
               hl_gto_l0stx            => c_tie_low,
               hl_gto_l1               => c_tie_low,
               hl_gto_l2               => c_tie_low,
               hl_gto_l0stxfts         => c_tie_low,
               hl_gto_lbk              => c_tie_low,
               hl_gto_rcvry            => c_tie_low,
               hl_gto_cfg              => c_tie_low,
               no_pcie_train           => c_tie_low,
               tx_dllp_val             => c_tie_low_byte(1 downto 0),
               tx_pmtype               => c_tie_low_byte(2 downto 0),
               tx_vsd_data             => c_tie_low_dword(23 downto 0),
               tx_req_vc0              => ix_tx_req,
               tx_data_vc0             => ix_tx_data,
               tx_st_vc0               => ix_tx_st,
               tx_end_vc0              => ix_tx_end,
               tx_nlfy_vc0             => c_tie_low,
               ph_buf_status_vc0       => c_tie_low,
               pd_buf_status_vc0       => c_tie_low,
               nph_buf_status_vc0      => c_tie_low,
               npd_buf_status_vc0      => c_tie_low,
               ph_processed_vc0        => ix_fc_processed_ph,
               pd_processed_vc0        => ix_fc_processed_pd,
               nph_processed_vc0       => ix_fc_processed_nph,
               npd_processed_vc0       => ix_fc_processed_npd,
               pd_num_vc0              => ix_fc_num_pd,
               npd_num_vc0             => ix_fc_num_npd,
               cmpln_tout              => c_tie_low,
               cmpltr_abort_np         => c_tie_low,
               cmpltr_abort_p          => c_tie_low,
               unexp_cmpln             => c_tie_low,
               ur_np_ext               => c_tie_low,
               ur_p_ext                => c_tie_low,
               np_req_pend             => c_tie_low,
               pme_status              => c_tie_low,
               tx_lbk_data             => c_tie_low_hword,
               tx_lbk_kcntl            => c_tie_low_byte(1 downto 0),
               
               tx_lbk_rdy              => open,
               rx_lbk_data             => open,
               rx_lbk_kcntl            => open,
               tx_dllp_sent            => open,
               rxdp_pmd_type           => open,
               rxdp_vsd_data           => open,
               rxdp_dllp_val           => open,
               phy_pol_compliance      => open,
               phy_ltssm_state         => ox_phy_ltssm_state,
               tx_rdy_vc0              => ox_tx_rdy,
               tx_ca_ph_vc0            => ox_tx_ca_ph,
               tx_ca_pd_vc0            => ox_tx_ca_pd,
               tx_ca_nph_vc0           => ox_tx_ca_nph,
               tx_ca_npd_vc0           => ox_tx_ca_npd,
               tx_ca_cplh_vc0          => ox_tx_ca_cplh,
               tx_ca_cpld_vc0          => ox_tx_ca_cpld,
               tx_ca_p_recheck_vc0     => ox_tx_ca_p_recheck,
               tx_ca_cpl_recheck_vc0   => ox_tx_ca_cpl_recheck,
               rx_data_vc0             => ox_rx_data,
               rx_st_vc0               => ox_rx_st,
               rx_end_vc0              => ox_rx_end,
               rx_us_req_vc0           => open,
               rx_malf_tlp_vc0         => open,
               rx_bar_hit              => ox_rx_bar_hit,
               mm_enable               => ox_mm_enable,
               msi_enable              => ox_msi_enable,
               bus_num                 => ox_bus_num,
               dev_num                 => ox_dev_num,
               func_num                => ox_func_num,
               pm_power_state          => open,
               pme_en                  => open,
               cmd_reg_out             => ox_cmd_reg_out,
               dev_cntl_out            => ox_dev_cntl_out,
               lnk_cntl_out            => ox_lnk_cntl_out,
               dl_inactive             => open,
               dl_init                 => open,
               dl_active               => open,
               dl_up                   => ox_dl_up,
               sys_clk_125             => ox_clk_125,
               sci_wrdata              => c_tie_low_byte,
               sci_addr                => c_tie_low_byte(5 downto 0),
               sci_wrn                 => c_tie_high,
               sci_en                  => c_tie_low,
               sci_sel                 => c_tie_low,
               sci_en_ch0              => c_tie_low,
               sci_sel_ch0             => c_tie_low,
               sci_rd                  => c_tie_low,
               sci_rddata              => open
               );  
      End Generate;
      
      U1_V5_X :
      if g_ip_rev_id = "V5_x" Generate     
         Component pcie_x1_top
               -- Component description of older PCIe Cores, Rev 5.x
               --
               -- Module generated by ipExpress. Component name must match ipExpress name
               -- There is normally no need to change the port declarations
               --
               -- Based on Lattice template file found at location <ip_dir>/pcie_eval/<ip_name>/src/top/<ip_name>_eval_top.v
            Port (
               refclkp                 : in std_logic;
               refclkn                 : in std_logic;
               rst_n                   : in std_logic;
               hdinp0                  : in std_logic;
               hdinn0                  : in std_logic;
               flip_lanes              : in std_logic;
               inta_n                  : in std_logic;
               msi                     : in std_logic_vector(7 downto 0);
               force_lsm_active        : in std_logic;
               force_rec_ei            : in std_logic;
               force_phy_status        : in std_logic;
               force_disable_scr       : in std_logic;
               hl_snd_beacon           : in std_logic;
               hl_disable_scr          : in std_logic;
               hl_gto_dis              : in std_logic;
               hl_gto_det              : in std_logic;
               hl_gto_hrst             : in std_logic;
               hl_gto_l0stx            : in std_logic;
               hl_gto_l1               : in std_logic;
               hl_gto_l2               : in std_logic;
               hl_gto_l0stxfts         : in std_logic;
               hl_gto_lbk              : in std_logic;
               hl_gto_rcvry            : in std_logic;
               hl_gto_cfg              : in std_logic;
               no_pcie_train           : in std_logic;
               tx_dllp_val             : in std_logic_vector(1 downto 0);
               tx_pmtype               : in std_logic_vector(2 downto 0);
               tx_vsd_data             : in std_logic_vector(23 downto 0);
               tx_req_vc0              : in std_logic;
               tx_data_vc0             : in std_logic_vector(15 downto 0);
               tx_st_vc0               : in std_logic;
               tx_end_vc0              : in std_logic;
               tx_nlfy_vc0             : in std_logic;
               ph_buf_status_vc0       : in std_logic;
               pd_buf_status_vc0       : in std_logic;
               nph_buf_status_vc0      : in std_logic;
               npd_buf_status_vc0      : in std_logic;
               ph_processed_vc0        : in std_logic;
               pd_processed_vc0        : in std_logic;
               nph_processed_vc0       : in std_logic;
               npd_processed_vc0       : in std_logic;
               pd_num_vc0              : in std_logic_vector(7 downto 0);
               npd_num_vc0             : in std_logic_vector(7 downto 0);
               cmpln_tout              : in std_logic;
               cmpltr_abort_np         : in std_logic;
               cmpltr_abort_p          : in std_logic;
               unexp_cmpln             : in std_logic;
               ur_np_ext               : in std_logic;
               ur_p_ext                : in std_logic;
               np_req_pend             : in std_logic;
               pme_status              : in std_logic;
               tx_lbk_data             : in std_logic_vector(15 downto 0);
               tx_lbk_kcntl            : in std_logic_vector(1 downto 0);

               hdoutp0                 : out std_logic;
               hdoutn0                 : out std_logic;
               tx_lbk_rdy              : out std_logic;
               rx_lbk_data             : out std_logic_vector(15 downto 0);
               rx_lbk_kcntl            : out std_logic_vector(1 downto 0);
               tx_dllp_sent            : out std_logic;
               rxdp_pmd_type           : out std_logic_vector(2 downto 0);
               rxdp_vsd_data           : out std_logic_vector(23 downto 0);
               rxdp_dllp_val           : out std_logic_vector(1 downto 0);
               phy_pol_compliance      : out std_logic;
               phy_ltssm_state         : out std_logic_vector(3 downto 0);
               phy_ltssm_substate      : out std_logic_vector(2 downto 0);
               tx_rdy_vc0              : out std_logic;
               tx_ca_ph_vc0            : out std_logic_vector(8 downto 0);
               tx_ca_pd_vc0            : out std_logic_vector(12 downto 0);
               tx_ca_nph_vc0           : out std_logic_vector(8 downto 0);
               tx_ca_npd_vc0           : out std_logic_vector(12 downto 0);
               tx_ca_cplh_vc0          : out std_logic_vector(8 downto 0);
               tx_ca_cpld_vc0          : out std_logic_vector(12 downto 0);
               tx_ca_p_recheck_vc0     : out std_logic;
               tx_ca_cpl_recheck_vc0   : out std_logic;
               rx_data_vc0             : out std_logic_vector(15 downto 0);
               rx_st_vc0               : out std_logic;
               rx_end_vc0              : out std_logic;
               rx_us_req_vc0           : out std_logic;
               rx_malf_tlp_vc0         : out std_logic;
               rx_bar_hit              : out std_logic_vector(6 downto 0);
               mm_enable               : out std_logic_vector(2 downto 0);
               msi_enable              : out std_logic;
               bus_num                 : out std_logic_vector(7 downto 0);
               dev_num                 : out std_logic_vector(4 downto 0);
               func_num                : out std_logic_vector(2 downto 0);
               pm_power_state          : out std_logic_vector(1 downto 0);
               pme_en                  : out std_logic;
               cmd_reg_out             : out std_logic_vector(5 downto 0);
               dev_cntl_out            : out std_logic_vector(14 downto 0);
               lnk_cntl_out            : out std_logic_vector(7 downto 0);
               dl_inactive             : out std_logic;
               dl_init                 : out std_logic;
               dl_active               : out std_logic;
               dl_up                   : out std_logic;
               irst_n                  : out std_logic;
               sys_clk_125             : out std_logic       
               );
         End Component;      
   Begin
         U1_PCIE:
         pcie_x1_top
            Port Map (
               refclkp                 => ix_refclkp,
               refclkn                 => ix_refclkn,
               rst_n                   => ix_rst_n,
               hdinp0                  => ix_hdinp0,
               hdinn0                  => ix_hdinn0,

               flip_lanes              => c_tie_low,
               inta_n                  => s_rtl_inta_n,
               msi                     => ix_msi_req,
               force_lsm_active        => c_tie_low,
               force_rec_ei            => c_tie_low,
               force_phy_status        => c_tie_low,
               force_disable_scr       => c_tie_low,
               hl_snd_beacon           => c_tie_low,
               hl_disable_scr          => c_tie_low,
               hl_gto_dis              => c_tie_low,
               hl_gto_det              => c_tie_low,
               hl_gto_hrst             => c_tie_low,
               hl_gto_l0stx            => c_tie_low,
               hl_gto_l1               => c_tie_low,
               hl_gto_l2               => c_tie_low,
               hl_gto_l0stxfts         => c_tie_low,
               hl_gto_lbk              => c_tie_low,
               hl_gto_rcvry            => c_tie_low,
               hl_gto_cfg              => c_tie_low,
               no_pcie_train           => c_tie_low,
               tx_dllp_val             => c_tie_low_byte(1 downto 0),
               tx_pmtype               => c_tie_low_byte(2 downto 0),
               tx_vsd_data             => c_tie_low_dword(23 downto 0),
               tx_req_vc0              => ix_tx_req,
               tx_data_vc0             => ix_tx_data,
               tx_st_vc0               => ix_tx_st,
               tx_end_vc0              => ix_tx_end,
               tx_nlfy_vc0             => c_tie_low,
               ph_buf_status_vc0       => c_tie_low,
               pd_buf_status_vc0       => c_tie_low,
               nph_buf_status_vc0      => c_tie_low,
               npd_buf_status_vc0      => c_tie_low,
               ph_processed_vc0        => ix_fc_processed_ph,
               pd_processed_vc0        => ix_fc_processed_pd,
               nph_processed_vc0       => ix_fc_processed_nph,
               npd_processed_vc0       => ix_fc_processed_npd,
               pd_num_vc0              => ix_fc_num_pd,
               npd_num_vc0             => ix_fc_num_npd,
               cmpln_tout              => c_tie_low,
               cmpltr_abort_np         => c_tie_low,
               cmpltr_abort_p          => c_tie_low,
               unexp_cmpln             => c_tie_low,
               ur_np_ext               => c_tie_low,
               ur_p_ext                => c_tie_low,
               np_req_pend             => c_tie_low,
               pme_status              => c_tie_low,
               tx_lbk_data             => c_tie_low_hword,
               tx_lbk_kcntl            => c_tie_low_byte(1 downto 0),

               hdoutp0                 => ox_hdoutp0,
               hdoutn0                 => ox_hdoutn0,
               tx_lbk_rdy              => open,
               rx_lbk_data             => open,
               rx_lbk_kcntl            => open,
               tx_dllp_sent            => open,
               rxdp_pmd_type           => open,
               rxdp_vsd_data           => open,
               rxdp_dllp_val           => open,
               phy_pol_compliance      => open,
               phy_ltssm_state         => ox_phy_ltssm_state,
               phy_ltssm_substate      => open,
               tx_rdy_vc0              => ox_tx_rdy,
               tx_ca_ph_vc0            => ox_tx_ca_ph,
               tx_ca_pd_vc0            => ox_tx_ca_pd,
               tx_ca_nph_vc0           => ox_tx_ca_nph,
               tx_ca_npd_vc0           => ox_tx_ca_npd,
               tx_ca_cplh_vc0          => ox_tx_ca_cplh,
               tx_ca_cpld_vc0          => ox_tx_ca_cpld,
               tx_ca_p_recheck_vc0     => ox_tx_ca_p_recheck,
               tx_ca_cpl_recheck_vc0   => ox_tx_ca_cpl_recheck,
               rx_data_vc0             => ox_rx_data,
               rx_st_vc0               => ox_rx_st,
               rx_end_vc0              => ox_rx_end,
               rx_us_req_vc0           => open,
               rx_malf_tlp_vc0         => open,
               rx_bar_hit              => ox_rx_bar_hit,
               mm_enable               => ox_mm_enable,
               msi_enable              => ox_msi_enable,
               bus_num                 => ox_bus_num,
               dev_num                 => ox_dev_num,
               func_num                => ox_func_num,
               pm_power_state          => open,
               pme_en                  => open,
               cmd_reg_out             => ox_cmd_reg_out,
               dev_cntl_out            => ox_dev_cntl_out,
               lnk_cntl_out            => ox_lnk_cntl_out,
               dl_inactive             => open,
               dl_init                 => open,
               dl_active               => open,
               dl_up                   => ox_dl_up,
               irst_n                  => open,
               sys_clk_125             => ox_clk_125
               );         
      End Generate;
   End Generate;
   
   U1_ECP5:
   if g_tech_lib = "ECP5UM" Generate
      
      U1_GEN1:
      if not g_pcie_gen2 Generate
         signal s_u1_refclk   : std_logic;
         
      begin
         U1_PCIE:            
         pcie_x1_e5
            Port Map (
               x_cref_refclkn                => ix_refclkn,
               x_cref_refclkp                => ix_refclkp,
               x_pcie_cmpln_tout             => c_tie_low,
               x_pcie_cmpltr_abort_np        => c_tie_low,
               x_pcie_cmpltr_abort_p         => c_tie_low,
               x_pcie_flip_lanes             => c_tie_low,
               x_pcie_force_disable_scr      => c_tie_low,
               x_pcie_force_lsm_active       => c_tie_low,
               x_pcie_force_phy_status       => c_tie_low,
               x_pcie_force_rec_ei           => c_tie_low,
               x_pcie_hdinn0                 => ix_hdinn0,
               x_pcie_hdinp0                 => ix_hdinp0,
               x_pcie_hl_disable_scr         => c_tie_low,
               x_pcie_hl_gto_cfg             => c_tie_low,
               x_pcie_hl_gto_det             => c_tie_low,
               x_pcie_hl_gto_dis             => c_tie_low,
               x_pcie_hl_gto_hrst            => c_tie_low,
               x_pcie_hl_gto_l0stx           => c_tie_low,
               x_pcie_hl_gto_l0stxfts        => c_tie_low,
               x_pcie_hl_gto_l1              => c_tie_low,
               x_pcie_hl_gto_l2              => c_tie_low,
               x_pcie_hl_gto_lbk             => c_tie_low,
               x_pcie_hl_gto_rcvry           => c_tie_low,
               x_pcie_hl_snd_beacon          => c_tie_low,
               x_pcie_inta_n                 => s_rtl_inta_n,
               x_pcie_msi                    => ix_msi_req,
               x_pcie_no_pcie_train          => c_tie_low,
               x_pcie_np_req_pend            => c_tie_low,
               x_pcie_npd_buf_status_vc0     => c_tie_low,
               x_pcie_npd_num_vc0            => ix_fc_num_npd,
               x_pcie_npd_processed_vc0      => ix_fc_processed_npd,
               x_pcie_nph_buf_status_vc0     => c_tie_low,
               x_pcie_nph_processed_vc0      => ix_fc_processed_nph,
               x_pcie_pd_buf_status_vc0      => c_tie_low,
               x_pcie_pd_num_vc0             => ix_fc_num_pd,
               x_pcie_pd_processed_vc0       => ix_fc_processed_pd,
               x_pcie_ph_buf_status_vc0      => c_tie_low,
               x_pcie_ph_processed_vc0       => ix_fc_processed_ph,
               x_pcie_pll_refclki            => s_u1_refclk,
               x_pcie_pme_status             => c_tie_low,
               x_pcie_rst_n                  => ix_rst_n,
               x_pcie_rxrefclk               => s_u1_refclk,
               x_pcie_sci_addr               => c_tie_low_byte(5 downto 0),
               x_pcie_sci_en                 => c_tie_low,
               x_pcie_sci_en_dual            => c_tie_low,
               x_pcie_sci_rd                 => c_tie_low,
               x_pcie_sci_sel                => c_tie_low,
               x_pcie_sci_sel_dual           => c_tie_low,
               x_pcie_sci_wrdata             => c_tie_low_byte,
               x_pcie_sci_wrn                => c_tie_high,
               x_pcie_tx_data_vc0            => ix_tx_data,
               x_pcie_tx_dllp_val            => c_tie_low_byte(1 downto 0),
               x_pcie_tx_end_vc0             => ix_tx_end,
               x_pcie_tx_lbk_data            => c_tie_low_hword,
               x_pcie_tx_lbk_kcntl           => c_tie_low_byte(1 downto 0),
               x_pcie_tx_nlfy_vc0            => c_tie_low,
               x_pcie_tx_pmtype              => c_tie_low_byte(2 downto 0),
               x_pcie_tx_req_vc0             => ix_tx_req,
               x_pcie_tx_st_vc0              => ix_tx_st,
               x_pcie_tx_vsd_data            => c_tie_low_dword(23 downto 0),
               x_pcie_unexp_cmpln            => c_tie_low,
               x_pcie_ur_np_ext              => c_tie_low,
               x_pcie_ur_p_ext               => c_tie_low,

               x_cref_refclko                => s_u1_refclk,
               x_pcie_bus_num                => ox_bus_num,
               x_pcie_cmd_reg_out            => ox_cmd_reg_out,
               x_pcie_dev_cntl_out           => ox_dev_cntl_out,
               x_pcie_dev_num                => ox_dev_num,
               x_pcie_dl_active              => open,
               x_pcie_dl_inactive            => open,
               x_pcie_dl_init                => open,
               x_pcie_dl_up                  => ox_dl_up,
               x_pcie_func_num               => ox_func_num,
               x_pcie_hdoutn0                => ox_hdoutn0,
               x_pcie_hdoutp0                => ox_hdoutp0,
               x_pcie_lnk_cntl_out           => ox_lnk_cntl_out,
               x_pcie_mm_enable              => ox_mm_enable,
               x_pcie_msi_enable             => ox_msi_enable,
               x_pcie_phy_ltssm_state        => ox_phy_ltssm_state,
               x_pcie_phy_pol_compliance     => open,
               x_pcie_pm_power_state         => open,
               x_pcie_pme_en                 => open,
               x_pcie_rx_bar_hit             => ox_rx_bar_hit,
               x_pcie_rx_data_vc0            => ox_rx_data,
               x_pcie_rx_end_vc0             => ox_rx_end,
               x_pcie_rx_lbk_data            => open,
               x_pcie_rx_lbk_kcntl           => open,
               x_pcie_rx_malf_tlp_vc0        => open,
               x_pcie_rx_st_vc0              => ox_rx_st,
               x_pcie_rx_us_req_vc0          => open,
               x_pcie_rxdp_dllp_val          => open,
               x_pcie_rxdp_pmd_type          => open,
               x_pcie_rxdp_vsd_data          => open,
               x_pcie_sci_int                => open,
               x_pcie_sci_rddata             => open,
               x_pcie_serdes_pdb             => open,
               x_pcie_serdes_rst_dual_c      => open,
               x_pcie_sys_clk_125            => ox_clk_125,
               x_pcie_tx_ca_cpl_recheck_vc0  => ox_tx_ca_cpl_recheck,
               x_pcie_tx_ca_cpld_vc0         => ox_tx_ca_cpld,
               x_pcie_tx_ca_cplh_vc0         => ox_tx_ca_cplh,
               x_pcie_tx_ca_npd_vc0          => ox_tx_ca_npd,
               x_pcie_tx_ca_nph_vc0          => ox_tx_ca_nph,
               x_pcie_tx_ca_p_recheck_vc0    => ox_tx_ca_p_recheck,
               x_pcie_tx_ca_pd_vc0           => ox_tx_ca_pd,
               x_pcie_tx_ca_ph_vc0           => ox_tx_ca_ph,
               x_pcie_tx_dllp_sent           => open,
               x_pcie_tx_lbk_rdy             => open,
               x_pcie_tx_pwrup_c             => open,
               x_pcie_tx_rdy_vc0             => ox_tx_rdy,
               x_pcie_tx_serdes_rst_c        => open
               );
      End Generate;

      U1_GEN2:
      if g_pcie_gen2 Generate
         signal s_u1_refclk   : std_logic;
      begin
         U1_PCIE:    
         pcie_x1_e5g2
            Port Map (
               x_cref_refclkn                => ix_refclkn,
               x_cref_refclkp                => ix_refclkp,
               x_pcie_cmpln_tout             => c_tie_low,
               x_pcie_cmpltr_abort_np        => c_tie_low,
               x_pcie_cmpltr_abort_p         => c_tie_low,
               x_pcie_flip_lanes             => c_tie_low,
               x_pcie_flr_rdy_in             => c_tie_low,
               x_pcie_force_disable_scr      => c_tie_low,
               x_pcie_force_lsm_active       => c_tie_low,
               x_pcie_force_phy_status       => c_tie_low,
               x_pcie_force_rec_ei           => c_tie_low,
               x_pcie_hdinn0                 => ix_hdinn0,
               x_pcie_hdinp0                 => ix_hdinp0,
               x_pcie_hl_disable_scr         => c_tie_low,
               x_pcie_hl_gto_cfg             => c_tie_low,
               x_pcie_hl_gto_det             => c_tie_low,
               x_pcie_hl_gto_dis             => c_tie_low,
               x_pcie_hl_gto_hrst            => c_tie_low,
               x_pcie_hl_gto_l0stx           => c_tie_low,
               x_pcie_hl_gto_l0stxfts        => c_tie_low,
               x_pcie_hl_gto_l1              => c_tie_low,
               x_pcie_hl_gto_l2              => c_tie_low,
               x_pcie_hl_gto_lbk             => c_tie_low_byte(1 downto 0),
               x_pcie_hl_gto_rcvry           => c_tie_low,
               x_pcie_hl_snd_beacon          => c_tie_low,
               x_pcie_inta_n                 => s_rtl_inta_n,
               x_pcie_msi                    => ix_msi_req,
               x_pcie_no_pcie_train          => c_tie_low,
               x_pcie_np_req_pend            => c_tie_low,
               x_pcie_npd_buf_status_vc0     => c_tie_low,
               x_pcie_npd_num_vc0            => ix_fc_num_npd,
               x_pcie_npd_processed_vc0      => ix_fc_processed_npd,
               x_pcie_nph_buf_status_vc0     => c_tie_low,
               x_pcie_nph_processed_vc0      => ix_fc_processed_nph,
               x_pcie_pd_buf_status_vc0      => c_tie_low,
               x_pcie_pd_num_vc0             => ix_fc_num_pd,
               x_pcie_pd_processed_vc0       => ix_fc_processed_pd,
               x_pcie_ph_buf_status_vc0      => c_tie_low,
               x_pcie_ph_processed_vc0       => ix_fc_processed_ph,
               x_pcie_pll_refclki            => s_u1_refclk,
               x_pcie_pme_status             => c_tie_low,
               x_pcie_rst_n                  => ix_rst_n,
               x_pcie_rxrefclk               => s_u1_refclk,
               x_pcie_tx_data_vc0            => c_tie_low_qword,  --ix_tx_data,
               x_pcie_tx_dllp_val            => c_tie_low_byte(1 downto 0),
               x_pcie_tx_dwen_vc0            => c_tie_low,
               x_pcie_tx_end_vc0             => ix_tx_end,
               x_pcie_tx_lbk_data            => c_tie_low_qword,
               x_pcie_tx_lbk_kcntl           => c_tie_low_byte,
               x_pcie_tx_nlfy_vc0            => c_tie_low,
               x_pcie_tx_pmtype              => c_tie_low_byte(2 downto 0),
               x_pcie_tx_req_vc0             => ix_tx_req,
               x_pcie_tx_st_vc0              => ix_tx_st,
               x_pcie_tx_vsd_data            => c_tie_low_dword(23 downto 0),
               x_pcie_unexp_cmpln            => c_tie_low,
               x_pcie_ur_np_ext              => c_tie_low,
               x_pcie_ur_p_ext               => c_tie_low,

               x_cref_refclko                => s_u1_refclk,
               x_pcie_bus_num                => ox_bus_num,
               x_pcie_cmd_reg_out            => ox_cmd_reg_out,
               x_pcie_dev_cntl_2_out         => open,
               x_pcie_dev_cntl_out           => ox_dev_cntl_out,
               x_pcie_dev_num                => ox_dev_num,
               x_pcie_dl_active              => open,
               x_pcie_dl_inactive            => open,
               x_pcie_dl_init                => open,
               x_pcie_dl_up                  => ox_dl_up,
               x_pcie_func_num               => ox_func_num,
               x_pcie_hdoutn0                => ox_hdoutn0,
               x_pcie_hdoutp0                => ox_hdoutp0,
               x_pcie_initiate_flr           => open,
               x_pcie_lnk_cntl_out           => ox_lnk_cntl_out,
               x_pcie_mm_enable              => ox_mm_enable,
               x_pcie_msi_enable             => ox_msi_enable,
               x_pcie_phy_cfgln              => open,
               x_pcie_phy_cfgln_sum          => open,
               x_pcie_phy_ltssm_state        => ox_phy_ltssm_state,
               x_pcie_phy_pol_compliance     => open,
               x_pcie_pm_power_state         => open,
               x_pcie_pme_en                 => open,
               x_pcie_rx_bar_hit             => ox_rx_bar_hit,
               x_pcie_rx_data_vc0            => open, --ox_rx_data,
               x_pcie_rx_end_vc0             => ox_rx_end,
               x_pcie_rx_lbk_data            => open,
               x_pcie_rx_lbk_kcntl           => open,
               x_pcie_rx_malf_tlp_vc0        => open,
               x_pcie_rx_st_vc0              => ox_rx_st,
               x_pcie_rx_us_req_vc0          => open,
               x_pcie_rxdp_dllp_val          => open,
               x_pcie_rxdp_pmd_type          => open,
               x_pcie_rxdp_vsd_data          => open,
               x_pcie_sys_clk_125            => ox_clk_125,
               x_pcie_tx_ca_cpl_recheck_vc0  => ox_tx_ca_cpl_recheck,
               x_pcie_tx_ca_cpld_vc0         => ox_tx_ca_cpld,
               x_pcie_tx_ca_cplh_vc0         => ox_tx_ca_cplh,
               x_pcie_tx_ca_npd_vc0          => ox_tx_ca_npd,
               x_pcie_tx_ca_nph_vc0          => ox_tx_ca_nph,
               x_pcie_tx_ca_p_recheck_vc0    => ox_tx_ca_p_recheck,
               x_pcie_tx_ca_pd_vc0           => ox_tx_ca_pd,
               x_pcie_tx_ca_ph_vc0           => ox_tx_ca_ph,
               x_pcie_tx_dllp_sent           => open,
               x_pcie_tx_lbk_rdy             => open,
               x_pcie_tx_rdy_vc0             => ox_tx_rdy
               );         
      End Generate;
   End Generate;
   
--    U2_RST_GEN:
--    tspc_rst_gen_yog4
--    Port Map (
--       i_clk       => s_u1_refclk,
--       i_trip_ev   => c_tie_low,
--       
--       o_rst_n     => s_u2_rst_n
--       );
End Rtl;
