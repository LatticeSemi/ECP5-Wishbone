
--    
--    Copyright Ingenieurbuero Gardiner, 2021
--       https://www.ib-gardiner.eu
--       techsupport@ib-gardiner.eu
--
--    All Rights Reserved
--   
--------------------------------------------------------------------------------
--
-- File ID    : $Id: config_ae53_ecp2m_v5-p.vhd 43 2021-11-18 17:41:37Z  $
-- Generated  : $LastChangedDate: 2021-11-18 18:41:37 +0100 (Thu, 18 Nov 2021) $
-- Revision   : $LastChangedRevision: 43 $
--
--------------------------------------------------------------------------------
--
-- Description : 
--
--------------------------------------------------------------------------------

Package core_ae53_config is
   constant c_pcie_gen2          : boolean := false;
   constant c_pcie_ip_rev_id     : string := "V5_x";
   constant c_tech_lib           : string := "ECP2M";
End core_ae53_config;
