Entity versa_ecp3_tb is
End versa_ecp3_tb;
